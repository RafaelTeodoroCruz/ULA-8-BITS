<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>10.7,-133.205,324.75,-293.763</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>63.5,-203.5</position>
<output>
<ID>OUT_0</ID>271 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2</ID>
<type>DD_KEYPAD_HEX</type>
<position>113.5,-168</position>
<output>
<ID>OUT_0</ID>5 </output>
<output>
<ID>OUT_1</ID>6 </output>
<output>
<ID>OUT_2</ID>7 </output>
<output>
<ID>OUT_3</ID>17 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>DD_KEYPAD_HEX</type>
<position>116,-187.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>2 </output>
<output>
<ID>OUT_2</ID>3 </output>
<output>
<ID>OUT_3</ID>4 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>174,-144</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_LABEL</type>
<position>62.5,-216</position>
<gparam>LABEL_TEXT FLAGS</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>BI_ROM_12x16</type>
<position>146.5,-168</position>
<input>
<ID>ADDRESS_0</ID>1 </input>
<input>
<ID>ADDRESS_1</ID>2 </input>
<input>
<ID>ADDRESS_10</ID>20 </input>
<input>
<ID>ADDRESS_11</ID>21 </input>
<input>
<ID>ADDRESS_2</ID>3 </input>
<input>
<ID>ADDRESS_3</ID>4 </input>
<input>
<ID>ADDRESS_4</ID>5 </input>
<input>
<ID>ADDRESS_5</ID>6 </input>
<input>
<ID>ADDRESS_6</ID>7 </input>
<input>
<ID>ADDRESS_7</ID>17 </input>
<input>
<ID>ADDRESS_8</ID>18 </input>
<input>
<ID>ADDRESS_9</ID>19 </input>
<output>
<ID>DATA_OUT_0</ID>22 </output>
<output>
<ID>DATA_OUT_1</ID>23 </output>
<output>
<ID>DATA_OUT_2</ID>24 </output>
<output>
<ID>DATA_OUT_3</ID>29 </output>
<output>
<ID>DATA_OUT_4</ID>38 </output>
<output>
<ID>DATA_OUT_5</ID>42 </output>
<output>
<ID>DATA_OUT_6</ID>43 </output>
<output>
<ID>DATA_OUT_7</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:1 1</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:3 3</lparam>
<lparam>Address:4 4</lparam>
<lparam>Address:5 5</lparam>
<lparam>Address:6 6</lparam>
<lparam>Address:7 7</lparam>
<lparam>Address:8 8</lparam>
<lparam>Address:9 9</lparam>
<lparam>Address:16 10</lparam>
<lparam>Address:17 11</lparam>
<lparam>Address:18 12</lparam>
<lparam>Address:19 13</lparam>
<lparam>Address:20 14</lparam>
<lparam>Address:21 15</lparam>
<lparam>Address:22 16</lparam>
<lparam>Address:23 17</lparam>
<lparam>Address:24 18</lparam>
<lparam>Address:25 19</lparam>
<lparam>Address:32 20</lparam>
<lparam>Address:33 21</lparam>
<lparam>Address:34 22</lparam>
<lparam>Address:35 23</lparam>
<lparam>Address:36 24</lparam>
<lparam>Address:37 25</lparam>
<lparam>Address:38 26</lparam>
<lparam>Address:39 27</lparam>
<lparam>Address:40 28</lparam>
<lparam>Address:41 29</lparam>
<lparam>Address:48 30</lparam>
<lparam>Address:49 31</lparam>
<lparam>Address:50 32</lparam>
<lparam>Address:51 33</lparam>
<lparam>Address:52 34</lparam>
<lparam>Address:53 35</lparam>
<lparam>Address:54 36</lparam>
<lparam>Address:55 37</lparam>
<lparam>Address:56 38</lparam>
<lparam>Address:57 39</lparam>
<lparam>Address:64 40</lparam>
<lparam>Address:65 41</lparam>
<lparam>Address:66 42</lparam>
<lparam>Address:67 43</lparam>
<lparam>Address:68 44</lparam>
<lparam>Address:69 45</lparam>
<lparam>Address:70 46</lparam>
<lparam>Address:71 47</lparam>
<lparam>Address:72 48</lparam>
<lparam>Address:73 49</lparam>
<lparam>Address:80 50</lparam>
<lparam>Address:81 51</lparam>
<lparam>Address:82 52</lparam>
<lparam>Address:83 53</lparam>
<lparam>Address:84 54</lparam>
<lparam>Address:85 55</lparam>
<lparam>Address:86 56</lparam>
<lparam>Address:87 57</lparam>
<lparam>Address:88 58</lparam>
<lparam>Address:89 59</lparam>
<lparam>Address:96 60</lparam>
<lparam>Address:97 61</lparam>
<lparam>Address:98 62</lparam>
<lparam>Address:99 63</lparam>
<lparam>Address:100 64</lparam>
<lparam>Address:101 65</lparam>
<lparam>Address:102 66</lparam>
<lparam>Address:103 67</lparam>
<lparam>Address:104 68</lparam>
<lparam>Address:105 69</lparam>
<lparam>Address:112 70</lparam>
<lparam>Address:113 71</lparam>
<lparam>Address:114 72</lparam>
<lparam>Address:115 73</lparam>
<lparam>Address:116 74</lparam>
<lparam>Address:117 75</lparam>
<lparam>Address:118 76</lparam>
<lparam>Address:119 77</lparam>
<lparam>Address:120 78</lparam>
<lparam>Address:121 79</lparam>
<lparam>Address:128 80</lparam>
<lparam>Address:129 81</lparam>
<lparam>Address:130 82</lparam>
<lparam>Address:131 83</lparam>
<lparam>Address:132 84</lparam>
<lparam>Address:133 85</lparam>
<lparam>Address:134 86</lparam>
<lparam>Address:135 87</lparam>
<lparam>Address:136 88</lparam>
<lparam>Address:137 89</lparam>
<lparam>Address:144 90</lparam>
<lparam>Address:145 91</lparam>
<lparam>Address:146 92</lparam>
<lparam>Address:147 93</lparam>
<lparam>Address:148 94</lparam>
<lparam>Address:149 95</lparam>
<lparam>Address:150 96</lparam>
<lparam>Address:151 97</lparam>
<lparam>Address:152 98</lparam>
<lparam>Address:153 99</lparam>
<lparam>Address:256 100</lparam>
<lparam>Address:257 101</lparam>
<lparam>Address:258 102</lparam>
<lparam>Address:259 103</lparam>
<lparam>Address:260 104</lparam>
<lparam>Address:261 105</lparam>
<lparam>Address:262 106</lparam>
<lparam>Address:263 107</lparam>
<lparam>Address:264 108</lparam>
<lparam>Address:265 109</lparam>
<lparam>Address:272 110</lparam>
<lparam>Address:273 111</lparam>
<lparam>Address:274 112</lparam>
<lparam>Address:275 113</lparam>
<lparam>Address:276 114</lparam>
<lparam>Address:277 115</lparam>
<lparam>Address:278 116</lparam>
<lparam>Address:279 117</lparam>
<lparam>Address:280 118</lparam>
<lparam>Address:281 119</lparam>
<lparam>Address:288 120</lparam>
<lparam>Address:289 121</lparam>
<lparam>Address:290 122</lparam>
<lparam>Address:291 123</lparam>
<lparam>Address:292 124</lparam>
<lparam>Address:293 125</lparam>
<lparam>Address:294 126</lparam>
<lparam>Address:295 127</lparam>
<lparam>Address:296 128</lparam>
<lparam>Address:297 129</lparam>
<lparam>Address:304 130</lparam>
<lparam>Address:305 131</lparam>
<lparam>Address:306 132</lparam>
<lparam>Address:307 133</lparam>
<lparam>Address:308 134</lparam>
<lparam>Address:309 135</lparam>
<lparam>Address:310 136</lparam>
<lparam>Address:311 137</lparam>
<lparam>Address:312 138</lparam>
<lparam>Address:313 139</lparam>
<lparam>Address:320 140</lparam>
<lparam>Address:321 141</lparam>
<lparam>Address:322 142</lparam>
<lparam>Address:323 143</lparam>
<lparam>Address:324 144</lparam>
<lparam>Address:325 145</lparam>
<lparam>Address:326 146</lparam>
<lparam>Address:327 147</lparam>
<lparam>Address:328 148</lparam>
<lparam>Address:329 149</lparam>
<lparam>Address:336 150</lparam>
<lparam>Address:337 151</lparam>
<lparam>Address:338 152</lparam>
<lparam>Address:339 153</lparam>
<lparam>Address:340 154</lparam>
<lparam>Address:341 155</lparam>
<lparam>Address:342 156</lparam>
<lparam>Address:343 157</lparam>
<lparam>Address:344 158</lparam>
<lparam>Address:345 159</lparam>
<lparam>Address:352 160</lparam>
<lparam>Address:353 161</lparam>
<lparam>Address:354 162</lparam>
<lparam>Address:355 163</lparam>
<lparam>Address:356 164</lparam>
<lparam>Address:357 165</lparam>
<lparam>Address:358 166</lparam>
<lparam>Address:359 167</lparam>
<lparam>Address:360 168</lparam>
<lparam>Address:361 169</lparam>
<lparam>Address:368 170</lparam>
<lparam>Address:369 171</lparam>
<lparam>Address:370 172</lparam>
<lparam>Address:371 173</lparam>
<lparam>Address:372 174</lparam>
<lparam>Address:373 175</lparam>
<lparam>Address:374 176</lparam>
<lparam>Address:375 177</lparam>
<lparam>Address:376 178</lparam>
<lparam>Address:377 179</lparam>
<lparam>Address:384 180</lparam>
<lparam>Address:385 181</lparam>
<lparam>Address:386 182</lparam>
<lparam>Address:387 183</lparam>
<lparam>Address:388 184</lparam>
<lparam>Address:389 185</lparam>
<lparam>Address:390 186</lparam>
<lparam>Address:391 187</lparam>
<lparam>Address:392 188</lparam>
<lparam>Address:393 189</lparam>
<lparam>Address:400 190</lparam>
<lparam>Address:401 191</lparam>
<lparam>Address:402 192</lparam>
<lparam>Address:403 193</lparam>
<lparam>Address:404 194</lparam>
<lparam>Address:405 195</lparam>
<lparam>Address:406 196</lparam>
<lparam>Address:407 197</lparam>
<lparam>Address:408 198</lparam>
<lparam>Address:409 199</lparam>
<lparam>Address:512 200</lparam>
<lparam>Address:513 201</lparam>
<lparam>Address:514 202</lparam>
<lparam>Address:515 203</lparam>
<lparam>Address:516 204</lparam>
<lparam>Address:517 205</lparam>
<lparam>Address:518 206</lparam>
<lparam>Address:519 207</lparam>
<lparam>Address:520 208</lparam>
<lparam>Address:521 209</lparam>
<lparam>Address:528 210</lparam>
<lparam>Address:529 211</lparam>
<lparam>Address:530 212</lparam>
<lparam>Address:531 213</lparam>
<lparam>Address:532 214</lparam>
<lparam>Address:533 215</lparam>
<lparam>Address:534 216</lparam>
<lparam>Address:535 217</lparam>
<lparam>Address:536 218</lparam>
<lparam>Address:537 219</lparam>
<lparam>Address:544 220</lparam>
<lparam>Address:545 221</lparam>
<lparam>Address:546 222</lparam>
<lparam>Address:547 223</lparam>
<lparam>Address:548 224</lparam>
<lparam>Address:549 225</lparam>
<lparam>Address:550 226</lparam>
<lparam>Address:551 227</lparam>
<lparam>Address:552 228</lparam>
<lparam>Address:553 229</lparam>
<lparam>Address:560 230</lparam>
<lparam>Address:561 231</lparam>
<lparam>Address:562 232</lparam>
<lparam>Address:563 233</lparam>
<lparam>Address:564 234</lparam>
<lparam>Address:565 235</lparam>
<lparam>Address:566 236</lparam>
<lparam>Address:567 237</lparam>
<lparam>Address:568 238</lparam>
<lparam>Address:569 239</lparam>
<lparam>Address:576 240</lparam>
<lparam>Address:577 241</lparam>
<lparam>Address:578 242</lparam>
<lparam>Address:579 243</lparam>
<lparam>Address:580 244</lparam>
<lparam>Address:581 245</lparam>
<lparam>Address:582 246</lparam>
<lparam>Address:583 247</lparam>
<lparam>Address:584 248</lparam>
<lparam>Address:585 249</lparam>
<lparam>Address:592 250</lparam>
<lparam>Address:593 251</lparam>
<lparam>Address:594 252</lparam>
<lparam>Address:595 253</lparam>
<lparam>Address:596 254</lparam>
<lparam>Address:597 255</lparam></gate>
<gate>
<ID>395</ID>
<type>DA_FROM</type>
<position>53,-235.5</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID v</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_DFF_LOW</type>
<position>195.5,-147</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUTINV_0</ID>11 </output>
<output>
<ID>OUT_0</ID>13 </output>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>396</ID>
<type>DA_FROM</type>
<position>53,-229</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID z</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>162,-144.5</position>
<gparam>LABEL_TEXT Push Button</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>397</ID>
<type>DA_FROM</type>
<position>53,-241.5</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID n</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND2</type>
<position>208,-145.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>398</ID>
<type>DA_FROM</type>
<position>53,-222</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c</lparam></gate>
<gate>
<ID>9</ID>
<type>DE_TO</type>
<position>215,-145</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID sinc</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>201.5,-142.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>11</ID>
<type>BB_CLOCK</type>
<position>180,-148</position>
<output>
<ID>CLK</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 10</lparam></gate>
<gate>
<ID>12</ID>
<type>DD_KEYPAD_HEX</type>
<position>116,-150.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<output>
<ID>OUT_1</ID>19 </output>
<output>
<ID>OUT_2</ID>20 </output>
<output>
<ID>OUT_3</ID>21 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>53,-192.5</position>
<gparam>LABEL_TEXT  G =X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1181</ID>
<type>DA_FROM</type>
<position>163.5,-247</position>
<input>
<ID>IN_0</ID>745 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID sinc</lparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>219.5,-153</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>1182</ID>
<type>DA_FROM</type>
<position>164,-265.5</position>
<input>
<ID>IN_0</ID>746 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>100,-164.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1185</ID>
<type>AA_LABEL</type>
<position>223.5,-195</position>
<gparam>LABEL_TEXT SAIDAS</gparam>
<gparam>TEXT_HEIGHT 7</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1186</ID>
<type>AA_LABEL</type>
<position>251,-227.5</position>
<gparam>LABEL_TEXT Display</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>68,-203.5</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1187</ID>
<type>AA_LABEL</type>
<position>242.5,-259</position>
<gparam>LABEL_TEXT LEDs em Binario</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>92.5,-203.5</position>
<output>
<ID>OUT_0</ID>269 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1188</ID>
<type>AA_LABEL</type>
<position>306,-283</position>
<gparam>LABEL_TEXT G1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>82.5,-203.5</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1189</ID>
<type>AA_AND2</type>
<position>298.5,-269.5</position>
<input>
<ID>IN_0</ID>748 </input>
<input>
<ID>IN_1</ID>758 </input>
<output>
<ID>OUT</ID>760 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>78,-203.5</position>
<output>
<ID>OUT_0</ID>270 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1190</ID>
<type>DA_FROM</type>
<position>290.5,-267.5</position>
<input>
<ID>IN_0</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g1</lparam></gate>
<gate>
<ID>1191</ID>
<type>DA_FROM</type>
<position>290.5,-271.5</position>
<input>
<ID>IN_0</ID>758 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>24</ID>
<type>DE_TO</type>
<position>97,-203.5</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1192</ID>
<type>GA_LED</type>
<position>302,-283.5</position>
<input>
<ID>N_in0</ID>760 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>57,-190</position>
<gparam>LABEL_TEXT G = X + 1 </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1193</ID>
<type>AA_LABEL</type>
<position>273,-283</position>
<gparam>LABEL_TEXT G3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1194</ID>
<type>AA_AND2</type>
<position>265.5,-269.5</position>
<input>
<ID>IN_0</ID>764 </input>
<input>
<ID>IN_1</ID>765 </input>
<output>
<ID>OUT</ID>766 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1195</ID>
<type>DA_FROM</type>
<position>257.5,-267.5</position>
<input>
<ID>IN_0</ID>764 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g3</lparam></gate>
<gate>
<ID>1196</ID>
<type>DA_FROM</type>
<position>257.5,-271.5</position>
<input>
<ID>IN_0</ID>765 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>1586</ID>
<type>AA_LABEL</type>
<position>247.5,-153.5</position>
<gparam>LABEL_TEXT GRUPO 7 </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1197</ID>
<type>GA_LED</type>
<position>269,-283.5</position>
<input>
<ID>N_in0</ID>766 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1198</ID>
<type>AA_LABEL</type>
<position>289.5,-283</position>
<gparam>LABEL_TEXT G2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1588</ID>
<type>AA_LABEL</type>
<position>279,-148</position>
<gparam>LABEL_TEXT ALGEBRA BOOLEANA E CIRCUITOS - G12 MATUTINO</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1199</ID>
<type>AA_AND2</type>
<position>282,-269.5</position>
<input>
<ID>IN_0</ID>761 </input>
<input>
<ID>IN_1</ID>762 </input>
<output>
<ID>OUT</ID>763 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>116,-142.5</position>
<gparam>LABEL_TEXT Centena</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1589</ID>
<type>AA_LABEL</type>
<position>275.5,-167</position>
<gparam>LABEL_TEXT Nome: Leonardo Aquino Cruz     RA:10445016 </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1200</ID>
<type>DA_FROM</type>
<position>274,-267.5</position>
<input>
<ID>IN_0</ID>761 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g2</lparam></gate>
<gate>
<ID>1590</ID>
<type>AA_LABEL</type>
<position>274,-171.5</position>
<gparam>LABEL_TEXT Nome: Rafael Teodoro Cruz     RA:10723258 </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1201</ID>
<type>DA_FROM</type>
<position>274,-271.5</position>
<input>
<ID>IN_0</ID>762 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>1591</ID>
<type>AA_LABEL</type>
<position>280,-176</position>
<gparam>LABEL_TEXT Nome: Joao Pedro Pereira Monteiro     RA:10727509 </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1202</ID>
<type>GA_LED</type>
<position>285.5,-283.5</position>
<input>
<ID>N_in0</ID>763 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>813</ID>
<type>GA_LED</type>
<position>61,-229</position>
<input>
<ID>N_in0</ID>494 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1592</ID>
<type>AA_LABEL</type>
<position>274.5,-180.5</position>
<gparam>LABEL_TEXT Nome: Joao Pedro Honorato     RA:10726497 </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1203</ID>
<type>AA_LABEL</type>
<position>239.5,-283</position>
<gparam>LABEL_TEXT G5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1593</ID>
<type>AA_LABEL</type>
<position>271.5,-160</position>
<gparam>LABEL_TEXT -Projeto 2 - ULA 8 BITS-</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1204</ID>
<type>AA_AND2</type>
<position>232,-269.5</position>
<input>
<ID>IN_0</ID>770 </input>
<input>
<ID>IN_1</ID>771 </input>
<output>
<ID>OUT</ID>772 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>815</ID>
<type>GA_LED</type>
<position>61,-241.5</position>
<input>
<ID>N_in0</ID>495 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1205</ID>
<type>DA_FROM</type>
<position>224,-267.5</position>
<input>
<ID>IN_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g5</lparam></gate>
<gate>
<ID>1206</ID>
<type>DA_FROM</type>
<position>224,-271.5</position>
<input>
<ID>IN_0</ID>771 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>817</ID>
<type>AA_LABEL</type>
<position>66,-228.5</position>
<gparam>LABEL_TEXT Zero</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>252.5,-241.5</position>
<input>
<ID>IN_0</ID>345 </input>
<input>
<ID>IN_1</ID>344 </input>
<input>
<ID>IN_2</ID>343 </input>
<input>
<ID>IN_3</ID>342 </input>
<input>
<ID>IN_4</ID>341 </input>
<input>
<ID>IN_5</ID>340 </input>
<input>
<ID>IN_6</ID>339 </input>
<input>
<ID>IN_7</ID>338 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1207</ID>
<type>GA_LED</type>
<position>235.5,-283.5</position>
<input>
<ID>N_in0</ID>772 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>429</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>233.5,-242.5</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>309 </input>
<input>
<ID>IN_2</ID>308 </input>
<input>
<ID>IN_3</ID>307 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1208</ID>
<type>AA_LABEL</type>
<position>256,-283</position>
<gparam>LABEL_TEXT G4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>819</ID>
<type>AA_LABEL</type>
<position>69.5,-241</position>
<gparam>LABEL_TEXT Negative</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1209</ID>
<type>AA_AND2</type>
<position>248.5,-269.5</position>
<input>
<ID>IN_0</ID>767 </input>
<input>
<ID>IN_1</ID>768 </input>
<output>
<ID>OUT</ID>769 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1210</ID>
<type>DA_FROM</type>
<position>240.5,-267.5</position>
<input>
<ID>IN_0</ID>767 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g4</lparam></gate>
<gate>
<ID>1211</ID>
<type>DA_FROM</type>
<position>240.5,-271.5</position>
<input>
<ID>IN_0</ID>768 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>1212</ID>
<type>GA_LED</type>
<position>252,-283.5</position>
<input>
<ID>N_in0</ID>769 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1213</ID>
<type>AA_LABEL</type>
<position>206.5,-283</position>
<gparam>LABEL_TEXT G7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1214</ID>
<type>AA_AND2</type>
<position>199,-269.5</position>
<input>
<ID>IN_0</ID>811 </input>
<input>
<ID>IN_1</ID>812 </input>
<output>
<ID>OUT</ID>813 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>DE_TO</type>
<position>176,-187.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>62</ID>
<type>DE_TO</type>
<position>176,-189.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>65</ID>
<type>DE_TO</type>
<position>176,-191.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>66</ID>
<type>DE_TO</type>
<position>176,-193.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>68</ID>
<type>DE_TO</type>
<position>176,-179.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>69</ID>
<type>DE_TO</type>
<position>176,-181.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>70</ID>
<type>DE_TO</type>
<position>176,-183.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>74</ID>
<type>DE_TO</type>
<position>176,-185.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>114,-160</position>
<gparam>LABEL_TEXT Dez</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>115.5,-179</position>
<gparam>LABEL_TEXT Unidade</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_TOGGLE</type>
<position>49,-203.5</position>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>89,-203</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>74.5,-203</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>AA_LABEL</type>
<position>60,-203</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>45.5,-203</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>AE_REGISTER8</type>
<position>165.5,-187</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>24 </input>
<input>
<ID>IN_3</ID>29 </input>
<input>
<ID>IN_4</ID>38 </input>
<input>
<ID>IN_5</ID>42 </input>
<input>
<ID>IN_6</ID>43 </input>
<input>
<ID>IN_7</ID>44 </input>
<output>
<ID>OUT_0</ID>8 </output>
<output>
<ID>OUT_1</ID>26 </output>
<output>
<ID>OUT_2</ID>25 </output>
<output>
<ID>OUT_3</ID>27 </output>
<output>
<ID>OUT_4</ID>28 </output>
<output>
<ID>OUT_5</ID>30 </output>
<output>
<ID>OUT_6</ID>31 </output>
<output>
<ID>OUT_7</ID>32 </output>
<input>
<ID>clock</ID>499 </input>
<input>
<ID>load</ID>484 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1309</ID>
<type>DA_FROM</type>
<position>191,-267.5</position>
<input>
<ID>IN_0</ID>811 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g7</lparam></gate>
<gate>
<ID>531</ID>
<type>GA_LED</type>
<position>61,-222</position>
<input>
<ID>N_in0</ID>489 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>532</ID>
<type>AA_LABEL</type>
<position>69.5,-221.5</position>
<gparam>LABEL_TEXT Carry-out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>536</ID>
<type>DA_FROM</type>
<position>162,-178</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID sinc</lparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>48,-159</position>
<input>
<ID>N_in0</ID>143 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1319</ID>
<type>DA_FROM</type>
<position>191,-271.5</position>
<input>
<ID>IN_0</ID>812 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>48,-156</position>
<input>
<ID>N_in0</ID>144 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1320</ID>
<type>GA_LED</type>
<position>202.5,-283.5</position>
<input>
<ID>N_in0</ID>813 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>GA_LED</type>
<position>48,-153</position>
<input>
<ID>N_in0</ID>145 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1321</ID>
<type>AA_LABEL</type>
<position>223,-283</position>
<gparam>LABEL_TEXT G6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>48,-162</position>
<input>
<ID>N_in0</ID>142 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1322</ID>
<type>AA_AND2</type>
<position>215.5,-269.5</position>
<input>
<ID>IN_0</ID>773 </input>
<input>
<ID>IN_1</ID>775 </input>
<output>
<ID>OUT</ID>810 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1323</ID>
<type>DA_FROM</type>
<position>207.5,-267.5</position>
<input>
<ID>IN_0</ID>773 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g6</lparam></gate>
<gate>
<ID>1324</ID>
<type>DA_FROM</type>
<position>207.5,-271.5</position>
<input>
<ID>IN_0</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>1325</ID>
<type>GA_LED</type>
<position>219,-283.5</position>
<input>
<ID>N_in0</ID>810 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>547</ID>
<type>AA_LABEL</type>
<position>322.5,-283</position>
<gparam>LABEL_TEXT G0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1327</ID>
<type>AA_LABEL</type>
<position>321,-288</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>BI_ROM_12x16</type>
<position>230.5,-218</position>
<input>
<ID>ADDRESS_0</ID>164 </input>
<input>
<ID>ADDRESS_1</ID>165 </input>
<input>
<ID>ADDRESS_2</ID>166 </input>
<input>
<ID>ADDRESS_3</ID>167 </input>
<input>
<ID>ADDRESS_4</ID>169 </input>
<input>
<ID>ADDRESS_5</ID>170 </input>
<input>
<ID>ADDRESS_6</ID>171 </input>
<input>
<ID>ADDRESS_7</ID>172 </input>
<output>
<ID>DATA_OUT_0</ID>345 </output>
<output>
<ID>DATA_OUT_1</ID>344 </output>
<output>
<ID>DATA_OUT_10</ID>308 </output>
<output>
<ID>DATA_OUT_11</ID>307 </output>
<output>
<ID>DATA_OUT_2</ID>343 </output>
<output>
<ID>DATA_OUT_3</ID>342 </output>
<output>
<ID>DATA_OUT_4</ID>341 </output>
<output>
<ID>DATA_OUT_5</ID>340 </output>
<output>
<ID>DATA_OUT_6</ID>339 </output>
<output>
<ID>DATA_OUT_7</ID>338 </output>
<output>
<ID>DATA_OUT_8</ID>310 </output>
<output>
<ID>DATA_OUT_9</ID>309 </output>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:1 1</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:3 3</lparam>
<lparam>Address:4 4</lparam>
<lparam>Address:5 5</lparam>
<lparam>Address:6 6</lparam>
<lparam>Address:7 7</lparam>
<lparam>Address:8 8</lparam>
<lparam>Address:9 9</lparam>
<lparam>Address:10 16</lparam>
<lparam>Address:11 17</lparam>
<lparam>Address:12 18</lparam>
<lparam>Address:13 19</lparam>
<lparam>Address:14 20</lparam>
<lparam>Address:15 21</lparam>
<lparam>Address:16 22</lparam>
<lparam>Address:17 23</lparam>
<lparam>Address:18 24</lparam>
<lparam>Address:19 25</lparam>
<lparam>Address:20 32</lparam>
<lparam>Address:21 33</lparam>
<lparam>Address:22 34</lparam>
<lparam>Address:23 35</lparam>
<lparam>Address:24 36</lparam>
<lparam>Address:25 37</lparam>
<lparam>Address:26 38</lparam>
<lparam>Address:27 39</lparam>
<lparam>Address:28 40</lparam>
<lparam>Address:29 41</lparam>
<lparam>Address:30 48</lparam>
<lparam>Address:31 49</lparam>
<lparam>Address:32 50</lparam>
<lparam>Address:33 51</lparam>
<lparam>Address:34 52</lparam>
<lparam>Address:35 53</lparam>
<lparam>Address:36 54</lparam>
<lparam>Address:37 55</lparam>
<lparam>Address:38 56</lparam>
<lparam>Address:39 57</lparam>
<lparam>Address:40 64</lparam>
<lparam>Address:41 65</lparam>
<lparam>Address:42 66</lparam>
<lparam>Address:43 67</lparam>
<lparam>Address:44 68</lparam>
<lparam>Address:45 69</lparam>
<lparam>Address:46 70</lparam>
<lparam>Address:47 71</lparam>
<lparam>Address:48 72</lparam>
<lparam>Address:49 73</lparam>
<lparam>Address:50 80</lparam>
<lparam>Address:51 81</lparam>
<lparam>Address:52 82</lparam>
<lparam>Address:53 83</lparam>
<lparam>Address:54 84</lparam>
<lparam>Address:55 85</lparam>
<lparam>Address:56 86</lparam>
<lparam>Address:57 87</lparam>
<lparam>Address:58 88</lparam>
<lparam>Address:59 89</lparam>
<lparam>Address:60 96</lparam>
<lparam>Address:61 97</lparam>
<lparam>Address:62 98</lparam>
<lparam>Address:63 99</lparam>
<lparam>Address:64 100</lparam>
<lparam>Address:65 101</lparam>
<lparam>Address:66 102</lparam>
<lparam>Address:67 103</lparam>
<lparam>Address:68 104</lparam>
<lparam>Address:69 105</lparam>
<lparam>Address:70 112</lparam>
<lparam>Address:71 113</lparam>
<lparam>Address:72 114</lparam>
<lparam>Address:73 115</lparam>
<lparam>Address:74 116</lparam>
<lparam>Address:75 117</lparam>
<lparam>Address:76 118</lparam>
<lparam>Address:77 119</lparam>
<lparam>Address:78 120</lparam>
<lparam>Address:79 121</lparam>
<lparam>Address:80 128</lparam>
<lparam>Address:81 129</lparam>
<lparam>Address:82 130</lparam>
<lparam>Address:83 131</lparam>
<lparam>Address:84 132</lparam>
<lparam>Address:85 133</lparam>
<lparam>Address:86 134</lparam>
<lparam>Address:87 135</lparam>
<lparam>Address:88 136</lparam>
<lparam>Address:89 137</lparam>
<lparam>Address:90 144</lparam>
<lparam>Address:91 145</lparam>
<lparam>Address:92 146</lparam>
<lparam>Address:93 147</lparam>
<lparam>Address:94 148</lparam>
<lparam>Address:95 149</lparam>
<lparam>Address:96 150</lparam>
<lparam>Address:97 151</lparam>
<lparam>Address:98 152</lparam>
<lparam>Address:99 153</lparam>
<lparam>Address:100 256</lparam>
<lparam>Address:101 257</lparam>
<lparam>Address:102 258</lparam>
<lparam>Address:103 259</lparam>
<lparam>Address:104 260</lparam>
<lparam>Address:105 261</lparam>
<lparam>Address:106 262</lparam>
<lparam>Address:107 263</lparam>
<lparam>Address:108 264</lparam>
<lparam>Address:109 265</lparam>
<lparam>Address:110 272</lparam>
<lparam>Address:111 273</lparam>
<lparam>Address:112 274</lparam>
<lparam>Address:113 275</lparam>
<lparam>Address:114 276</lparam>
<lparam>Address:115 277</lparam>
<lparam>Address:116 278</lparam>
<lparam>Address:117 279</lparam>
<lparam>Address:118 280</lparam>
<lparam>Address:119 281</lparam>
<lparam>Address:120 288</lparam>
<lparam>Address:121 289</lparam>
<lparam>Address:122 290</lparam>
<lparam>Address:123 291</lparam>
<lparam>Address:124 292</lparam>
<lparam>Address:125 293</lparam>
<lparam>Address:126 294</lparam>
<lparam>Address:127 295</lparam>
<lparam>Address:128 296</lparam>
<lparam>Address:129 297</lparam>
<lparam>Address:130 304</lparam>
<lparam>Address:131 305</lparam>
<lparam>Address:132 306</lparam>
<lparam>Address:133 307</lparam>
<lparam>Address:134 308</lparam>
<lparam>Address:135 309</lparam>
<lparam>Address:136 310</lparam>
<lparam>Address:137 311</lparam>
<lparam>Address:138 312</lparam>
<lparam>Address:139 313</lparam>
<lparam>Address:140 320</lparam>
<lparam>Address:141 321</lparam>
<lparam>Address:142 322</lparam>
<lparam>Address:143 323</lparam>
<lparam>Address:144 324</lparam>
<lparam>Address:145 325</lparam>
<lparam>Address:146 326</lparam>
<lparam>Address:147 327</lparam>
<lparam>Address:148 328</lparam>
<lparam>Address:149 329</lparam>
<lparam>Address:150 336</lparam>
<lparam>Address:151 337</lparam>
<lparam>Address:152 338</lparam>
<lparam>Address:153 339</lparam>
<lparam>Address:154 340</lparam>
<lparam>Address:155 341</lparam>
<lparam>Address:156 342</lparam>
<lparam>Address:157 343</lparam>
<lparam>Address:158 344</lparam>
<lparam>Address:159 345</lparam>
<lparam>Address:160 352</lparam>
<lparam>Address:161 353</lparam>
<lparam>Address:162 354</lparam>
<lparam>Address:163 355</lparam>
<lparam>Address:164 356</lparam>
<lparam>Address:165 357</lparam>
<lparam>Address:166 358</lparam>
<lparam>Address:167 359</lparam>
<lparam>Address:168 360</lparam>
<lparam>Address:169 361</lparam>
<lparam>Address:170 368</lparam>
<lparam>Address:171 369</lparam>
<lparam>Address:172 370</lparam>
<lparam>Address:173 371</lparam>
<lparam>Address:174 372</lparam>
<lparam>Address:175 373</lparam>
<lparam>Address:176 374</lparam>
<lparam>Address:177 375</lparam>
<lparam>Address:178 376</lparam>
<lparam>Address:179 377</lparam>
<lparam>Address:180 384</lparam>
<lparam>Address:181 385</lparam>
<lparam>Address:182 386</lparam>
<lparam>Address:183 387</lparam>
<lparam>Address:184 388</lparam>
<lparam>Address:185 389</lparam>
<lparam>Address:186 390</lparam>
<lparam>Address:187 391</lparam>
<lparam>Address:188 392</lparam>
<lparam>Address:189 393</lparam>
<lparam>Address:190 400</lparam>
<lparam>Address:191 401</lparam>
<lparam>Address:192 402</lparam>
<lparam>Address:193 403</lparam>
<lparam>Address:194 404</lparam>
<lparam>Address:195 405</lparam>
<lparam>Address:196 406</lparam>
<lparam>Address:197 407</lparam>
<lparam>Address:198 408</lparam>
<lparam>Address:199 409</lparam>
<lparam>Address:200 512</lparam>
<lparam>Address:201 513</lparam>
<lparam>Address:202 514</lparam>
<lparam>Address:203 515</lparam>
<lparam>Address:204 516</lparam>
<lparam>Address:205 517</lparam>
<lparam>Address:206 518</lparam>
<lparam>Address:207 519</lparam>
<lparam>Address:208 520</lparam>
<lparam>Address:209 521</lparam>
<lparam>Address:210 528</lparam>
<lparam>Address:211 529</lparam>
<lparam>Address:212 530</lparam>
<lparam>Address:213 531</lparam>
<lparam>Address:214 532</lparam>
<lparam>Address:215 533</lparam>
<lparam>Address:216 534</lparam>
<lparam>Address:217 535</lparam>
<lparam>Address:218 536</lparam>
<lparam>Address:219 537</lparam>
<lparam>Address:220 544</lparam>
<lparam>Address:221 545</lparam>
<lparam>Address:222 546</lparam>
<lparam>Address:223 547</lparam>
<lparam>Address:224 548</lparam>
<lparam>Address:225 549</lparam>
<lparam>Address:226 550</lparam>
<lparam>Address:227 551</lparam>
<lparam>Address:228 552</lparam>
<lparam>Address:229 553</lparam>
<lparam>Address:230 560</lparam>
<lparam>Address:231 561</lparam>
<lparam>Address:232 562</lparam>
<lparam>Address:233 563</lparam>
<lparam>Address:234 564</lparam>
<lparam>Address:235 565</lparam>
<lparam>Address:236 566</lparam>
<lparam>Address:237 567</lparam>
<lparam>Address:238 568</lparam>
<lparam>Address:239 569</lparam>
<lparam>Address:240 576</lparam>
<lparam>Address:241 577</lparam>
<lparam>Address:242 578</lparam>
<lparam>Address:243 579</lparam>
<lparam>Address:244 580</lparam>
<lparam>Address:245 581</lparam>
<lparam>Address:246 582</lparam>
<lparam>Address:247 583</lparam>
<lparam>Address:248 584</lparam>
<lparam>Address:249 585</lparam>
<lparam>Address:250 592</lparam>
<lparam>Address:251 593</lparam>
<lparam>Address:252 594</lparam>
<lparam>Address:253 595</lparam>
<lparam>Address:254 596</lparam>
<lparam>Address:255 597</lparam></gate>
<gate>
<ID>1328</ID>
<type>AA_LABEL</type>
<position>304.5,-288</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1329</ID>
<type>AA_LABEL</type>
<position>288,-288</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1330</ID>
<type>AA_LABEL</type>
<position>271.5,-288</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1331</ID>
<type>AA_LABEL</type>
<position>254.5,-288</position>
<gparam>LABEL_TEXT 16</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1332</ID>
<type>AA_LABEL</type>
<position>238,-288</position>
<gparam>LABEL_TEXT 32</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1333</ID>
<type>AA_LABEL</type>
<position>221.5,-288</position>
<gparam>LABEL_TEXT 64</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1334</ID>
<type>AA_LABEL</type>
<position>205,-288</position>
<gparam>LABEL_TEXT 128</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>AE_REGISTER8</type>
<position>212,-220.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>155 </input>
<input>
<ID>IN_2</ID>156 </input>
<input>
<ID>IN_3</ID>157 </input>
<input>
<ID>IN_4</ID>158 </input>
<input>
<ID>IN_5</ID>159 </input>
<input>
<ID>IN_6</ID>160 </input>
<input>
<ID>IN_7</ID>161 </input>
<output>
<ID>OUT_0</ID>164 </output>
<output>
<ID>OUT_1</ID>165 </output>
<output>
<ID>OUT_2</ID>166 </output>
<output>
<ID>OUT_3</ID>167 </output>
<output>
<ID>OUT_4</ID>169 </output>
<output>
<ID>OUT_5</ID>170 </output>
<output>
<ID>OUT_6</ID>171 </output>
<output>
<ID>OUT_7</ID>172 </output>
<input>
<ID>clock</ID>162 </input>
<input>
<ID>load</ID>163 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>170</ID>
<type>DA_FROM</type>
<position>196,-227</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g0</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>196,-225</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g1</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>196,-221</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g3</lparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>196,-217</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g5</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>196,-219</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g4</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>196,-223</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g2</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>196,-215</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g6</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>196,-213</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g7</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>209,-230</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>179</ID>
<type>EE_VDD</type>
<position>211,-211.5</position>
<output>
<ID>OUT_0</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>22.5,-189</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AA_LABEL</type>
<position>22.5,-192.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>AA_LABEL</type>
<position>22.5,-196</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>AA_LABEL</type>
<position>22.5,-199.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>AA_LABEL</type>
<position>22.5,-203</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>AA_LABEL</type>
<position>22.5,-206.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>22.5,-210</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>22.5,-213.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>22.5,-217</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>22.5,-220.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>22.5,-224</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>22.5,-227.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>22.5,-231</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>22.5,-234.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>22.5,-238</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>22.5,-241.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>607</ID>
<type>GA_LED</type>
<position>61,-235.5</position>
<input>
<ID>N_in0</ID>496 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>608</ID>
<type>AA_LABEL</type>
<position>69.5,-235</position>
<gparam>LABEL_TEXT Overflow</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>26,-189</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>26,-192.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_LABEL</type>
<position>26,-196</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>26,-199.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_LABEL</type>
<position>26,-217</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>224</ID>
<type>AA_LABEL</type>
<position>26,-220.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>AA_LABEL</type>
<position>26,-224</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>56,-187.5</position>
<gparam>LABEL_TEXT G = X - 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>DE_TO</type>
<position>53.5,-203.5</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_LABEL</type>
<position>56.5,-185</position>
<gparam>LABEL_TEXT  G = X + Y </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>229</ID>
<type>AA_LABEL</type>
<position>26,-227.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>230</ID>
<type>AA_LABEL</type>
<position>26,-203</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>26,-206.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_LABEL</type>
<position>26,-210</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>233</ID>
<type>AA_LABEL</type>
<position>26,-213.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>54,-182.5</position>
<gparam>LABEL_TEXT G = Y </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>235</ID>
<type>AA_LABEL</type>
<position>26,-231</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_LABEL</type>
<position>26,-234.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>237</ID>
<type>AA_LABEL</type>
<position>26,-238</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>238</ID>
<type>AA_LABEL</type>
<position>26,-241.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>239</ID>
<type>AA_LABEL</type>
<position>29.5,-189</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>240</ID>
<type>AA_LABEL</type>
<position>29.5,-192.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>29.5,-203</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>AA_LABEL</type>
<position>29.5,-206.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>AA_LABEL</type>
<position>29.5,-217</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>AA_LABEL</type>
<position>29.5,-220.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_LABEL</type>
<position>29.5,-231</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>635</ID>
<type>AA_LABEL</type>
<position>50,-140</position>
<gparam>LABEL_TEXT ULA</gparam>
<gparam>TEXT_HEIGHT 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>29.5,-234.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>AA_LABEL</type>
<position>56.5,-180</position>
<gparam>LABEL_TEXT G = Y + 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>AA_LABEL</type>
<position>55.5,-177.5</position>
<gparam>LABEL_TEXT  G= Y - 1 </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>GA_LED</type>
<position>48,-193</position>
<input>
<ID>N_in0</ID>286 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>60,-175</position>
<gparam>LABEL_TEXT G = X + Y' + 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>69.5,-152.5</position>
<gparam>LABEL_TEXT G = (X == Y) ? 0xFF : 0x00</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>GA_LED</type>
<position>48,-183</position>
<input>
<ID>N_in0</ID>318 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1033</ID>
<type>AA_LABEL</type>
<position>33,-189</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>255</ID>
<type>GA_LED</type>
<position>48,-180.5</position>
<input>
<ID>N_in0</ID>319 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1034</ID>
<type>DD_KEYPAD_HEX</type>
<position>115,-237</position>
<output>
<ID>OUT_0</ID>721 </output>
<output>
<ID>OUT_1</ID>722 </output>
<output>
<ID>OUT_2</ID>723 </output>
<output>
<ID>OUT_3</ID>725 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_LABEL</type>
<position>29.5,-196</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1035</ID>
<type>DD_KEYPAD_HEX</type>
<position>117.5,-256.5</position>
<output>
<ID>OUT_0</ID>689 </output>
<output>
<ID>OUT_1</ID>690 </output>
<output>
<ID>OUT_2</ID>719 </output>
<output>
<ID>OUT_3</ID>720 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_LABEL</type>
<position>29.5,-199.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1036</ID>
<type>BI_ROM_12x16</type>
<position>148,-237</position>
<input>
<ID>ADDRESS_0</ID>689 </input>
<input>
<ID>ADDRESS_1</ID>690 </input>
<input>
<ID>ADDRESS_10</ID>728 </input>
<input>
<ID>ADDRESS_11</ID>729 </input>
<input>
<ID>ADDRESS_2</ID>719 </input>
<input>
<ID>ADDRESS_3</ID>720 </input>
<input>
<ID>ADDRESS_4</ID>721 </input>
<input>
<ID>ADDRESS_5</ID>722 </input>
<input>
<ID>ADDRESS_6</ID>723 </input>
<input>
<ID>ADDRESS_7</ID>725 </input>
<input>
<ID>ADDRESS_8</ID>726 </input>
<input>
<ID>ADDRESS_9</ID>727 </input>
<output>
<ID>DATA_OUT_0</ID>730 </output>
<output>
<ID>DATA_OUT_1</ID>731 </output>
<output>
<ID>DATA_OUT_2</ID>732 </output>
<output>
<ID>DATA_OUT_3</ID>737 </output>
<output>
<ID>DATA_OUT_4</ID>741 </output>
<output>
<ID>DATA_OUT_5</ID>742 </output>
<output>
<ID>DATA_OUT_6</ID>743 </output>
<output>
<ID>DATA_OUT_7</ID>744 </output>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:1 1</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:3 3</lparam>
<lparam>Address:4 4</lparam>
<lparam>Address:5 5</lparam>
<lparam>Address:6 6</lparam>
<lparam>Address:7 7</lparam>
<lparam>Address:8 8</lparam>
<lparam>Address:9 9</lparam>
<lparam>Address:16 10</lparam>
<lparam>Address:17 11</lparam>
<lparam>Address:18 12</lparam>
<lparam>Address:19 13</lparam>
<lparam>Address:20 14</lparam>
<lparam>Address:21 15</lparam>
<lparam>Address:22 16</lparam>
<lparam>Address:23 17</lparam>
<lparam>Address:24 18</lparam>
<lparam>Address:25 19</lparam>
<lparam>Address:32 20</lparam>
<lparam>Address:33 21</lparam>
<lparam>Address:34 22</lparam>
<lparam>Address:35 23</lparam>
<lparam>Address:36 24</lparam>
<lparam>Address:37 25</lparam>
<lparam>Address:38 26</lparam>
<lparam>Address:39 27</lparam>
<lparam>Address:40 28</lparam>
<lparam>Address:41 29</lparam>
<lparam>Address:48 30</lparam>
<lparam>Address:49 31</lparam>
<lparam>Address:50 32</lparam>
<lparam>Address:51 33</lparam>
<lparam>Address:52 34</lparam>
<lparam>Address:53 35</lparam>
<lparam>Address:54 36</lparam>
<lparam>Address:55 37</lparam>
<lparam>Address:56 38</lparam>
<lparam>Address:57 39</lparam>
<lparam>Address:64 40</lparam>
<lparam>Address:65 41</lparam>
<lparam>Address:66 42</lparam>
<lparam>Address:67 43</lparam>
<lparam>Address:68 44</lparam>
<lparam>Address:69 45</lparam>
<lparam>Address:70 46</lparam>
<lparam>Address:71 47</lparam>
<lparam>Address:72 48</lparam>
<lparam>Address:73 49</lparam>
<lparam>Address:80 50</lparam>
<lparam>Address:81 51</lparam>
<lparam>Address:82 52</lparam>
<lparam>Address:83 53</lparam>
<lparam>Address:84 54</lparam>
<lparam>Address:85 55</lparam>
<lparam>Address:86 56</lparam>
<lparam>Address:87 57</lparam>
<lparam>Address:88 58</lparam>
<lparam>Address:89 59</lparam>
<lparam>Address:96 60</lparam>
<lparam>Address:97 61</lparam>
<lparam>Address:98 62</lparam>
<lparam>Address:99 63</lparam>
<lparam>Address:100 64</lparam>
<lparam>Address:101 65</lparam>
<lparam>Address:102 66</lparam>
<lparam>Address:103 67</lparam>
<lparam>Address:104 68</lparam>
<lparam>Address:105 69</lparam>
<lparam>Address:112 70</lparam>
<lparam>Address:113 71</lparam>
<lparam>Address:114 72</lparam>
<lparam>Address:115 73</lparam>
<lparam>Address:116 74</lparam>
<lparam>Address:117 75</lparam>
<lparam>Address:118 76</lparam>
<lparam>Address:119 77</lparam>
<lparam>Address:120 78</lparam>
<lparam>Address:121 79</lparam>
<lparam>Address:128 80</lparam>
<lparam>Address:129 81</lparam>
<lparam>Address:130 82</lparam>
<lparam>Address:131 83</lparam>
<lparam>Address:132 84</lparam>
<lparam>Address:133 85</lparam>
<lparam>Address:134 86</lparam>
<lparam>Address:135 87</lparam>
<lparam>Address:136 88</lparam>
<lparam>Address:137 89</lparam>
<lparam>Address:144 90</lparam>
<lparam>Address:145 91</lparam>
<lparam>Address:146 92</lparam>
<lparam>Address:147 93</lparam>
<lparam>Address:148 94</lparam>
<lparam>Address:149 95</lparam>
<lparam>Address:150 96</lparam>
<lparam>Address:151 97</lparam>
<lparam>Address:152 98</lparam>
<lparam>Address:153 99</lparam>
<lparam>Address:256 100</lparam>
<lparam>Address:257 101</lparam>
<lparam>Address:258 102</lparam>
<lparam>Address:259 103</lparam>
<lparam>Address:260 104</lparam>
<lparam>Address:261 105</lparam>
<lparam>Address:262 106</lparam>
<lparam>Address:263 107</lparam>
<lparam>Address:264 108</lparam>
<lparam>Address:265 109</lparam>
<lparam>Address:272 110</lparam>
<lparam>Address:273 111</lparam>
<lparam>Address:274 112</lparam>
<lparam>Address:275 113</lparam>
<lparam>Address:276 114</lparam>
<lparam>Address:277 115</lparam>
<lparam>Address:278 116</lparam>
<lparam>Address:279 117</lparam>
<lparam>Address:280 118</lparam>
<lparam>Address:281 119</lparam>
<lparam>Address:288 120</lparam>
<lparam>Address:289 121</lparam>
<lparam>Address:290 122</lparam>
<lparam>Address:291 123</lparam>
<lparam>Address:292 124</lparam>
<lparam>Address:293 125</lparam>
<lparam>Address:294 126</lparam>
<lparam>Address:295 127</lparam>
<lparam>Address:296 128</lparam>
<lparam>Address:297 129</lparam>
<lparam>Address:304 130</lparam>
<lparam>Address:305 131</lparam>
<lparam>Address:306 132</lparam>
<lparam>Address:307 133</lparam>
<lparam>Address:308 134</lparam>
<lparam>Address:309 135</lparam>
<lparam>Address:310 136</lparam>
<lparam>Address:311 137</lparam>
<lparam>Address:312 138</lparam>
<lparam>Address:313 139</lparam>
<lparam>Address:320 140</lparam>
<lparam>Address:321 141</lparam>
<lparam>Address:322 142</lparam>
<lparam>Address:323 143</lparam>
<lparam>Address:324 144</lparam>
<lparam>Address:325 145</lparam>
<lparam>Address:326 146</lparam>
<lparam>Address:327 147</lparam>
<lparam>Address:328 148</lparam>
<lparam>Address:329 149</lparam>
<lparam>Address:336 150</lparam>
<lparam>Address:337 151</lparam>
<lparam>Address:338 152</lparam>
<lparam>Address:339 153</lparam>
<lparam>Address:340 154</lparam>
<lparam>Address:341 155</lparam>
<lparam>Address:342 156</lparam>
<lparam>Address:343 157</lparam>
<lparam>Address:344 158</lparam>
<lparam>Address:345 159</lparam>
<lparam>Address:352 160</lparam>
<lparam>Address:353 161</lparam>
<lparam>Address:354 162</lparam>
<lparam>Address:355 163</lparam>
<lparam>Address:356 164</lparam>
<lparam>Address:357 165</lparam>
<lparam>Address:358 166</lparam>
<lparam>Address:359 167</lparam>
<lparam>Address:360 168</lparam>
<lparam>Address:361 169</lparam>
<lparam>Address:368 170</lparam>
<lparam>Address:369 171</lparam>
<lparam>Address:370 172</lparam>
<lparam>Address:371 173</lparam>
<lparam>Address:372 174</lparam>
<lparam>Address:373 175</lparam>
<lparam>Address:374 176</lparam>
<lparam>Address:375 177</lparam>
<lparam>Address:376 178</lparam>
<lparam>Address:377 179</lparam>
<lparam>Address:384 180</lparam>
<lparam>Address:385 181</lparam>
<lparam>Address:386 182</lparam>
<lparam>Address:387 183</lparam>
<lparam>Address:388 184</lparam>
<lparam>Address:389 185</lparam>
<lparam>Address:390 186</lparam>
<lparam>Address:391 187</lparam>
<lparam>Address:392 188</lparam>
<lparam>Address:393 189</lparam>
<lparam>Address:400 190</lparam>
<lparam>Address:401 191</lparam>
<lparam>Address:402 192</lparam>
<lparam>Address:403 193</lparam>
<lparam>Address:404 194</lparam>
<lparam>Address:405 195</lparam>
<lparam>Address:406 196</lparam>
<lparam>Address:407 197</lparam>
<lparam>Address:408 198</lparam>
<lparam>Address:409 199</lparam>
<lparam>Address:512 200</lparam>
<lparam>Address:513 201</lparam>
<lparam>Address:514 202</lparam>
<lparam>Address:515 203</lparam>
<lparam>Address:516 204</lparam>
<lparam>Address:517 205</lparam>
<lparam>Address:518 206</lparam>
<lparam>Address:519 207</lparam>
<lparam>Address:520 208</lparam>
<lparam>Address:521 209</lparam>
<lparam>Address:528 210</lparam>
<lparam>Address:529 211</lparam>
<lparam>Address:530 212</lparam>
<lparam>Address:531 213</lparam>
<lparam>Address:532 214</lparam>
<lparam>Address:533 215</lparam>
<lparam>Address:534 216</lparam>
<lparam>Address:535 217</lparam>
<lparam>Address:536 218</lparam>
<lparam>Address:537 219</lparam>
<lparam>Address:544 220</lparam>
<lparam>Address:545 221</lparam>
<lparam>Address:546 222</lparam>
<lparam>Address:547 223</lparam>
<lparam>Address:548 224</lparam>
<lparam>Address:549 225</lparam>
<lparam>Address:550 226</lparam>
<lparam>Address:551 227</lparam>
<lparam>Address:552 228</lparam>
<lparam>Address:553 229</lparam>
<lparam>Address:560 230</lparam>
<lparam>Address:561 231</lparam>
<lparam>Address:562 232</lparam>
<lparam>Address:563 233</lparam>
<lparam>Address:564 234</lparam>
<lparam>Address:565 235</lparam>
<lparam>Address:566 236</lparam>
<lparam>Address:567 237</lparam>
<lparam>Address:568 238</lparam>
<lparam>Address:569 239</lparam>
<lparam>Address:576 240</lparam>
<lparam>Address:577 241</lparam>
<lparam>Address:578 242</lparam>
<lparam>Address:579 243</lparam>
<lparam>Address:580 244</lparam>
<lparam>Address:581 245</lparam>
<lparam>Address:582 246</lparam>
<lparam>Address:583 247</lparam>
<lparam>Address:584 248</lparam>
<lparam>Address:585 249</lparam>
<lparam>Address:592 250</lparam>
<lparam>Address:593 251</lparam>
<lparam>Address:594 252</lparam>
<lparam>Address:595 253</lparam>
<lparam>Address:596 254</lparam>
<lparam>Address:597 255</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_LABEL</type>
<position>29.5,-210</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1037</ID>
<type>DD_KEYPAD_HEX</type>
<position>117.5,-219.5</position>
<output>
<ID>OUT_0</ID>726 </output>
<output>
<ID>OUT_1</ID>727 </output>
<output>
<ID>OUT_2</ID>728 </output>
<output>
<ID>OUT_3</ID>729 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_LABEL</type>
<position>29.5,-213.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1038</ID>
<type>AA_LABEL</type>
<position>101.5,-233.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>29.5,-224</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1039</ID>
<type>AA_LABEL</type>
<position>117.5,-211.5</position>
<gparam>LABEL_TEXT Centena</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AA_LABEL</type>
<position>29.5,-227.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1040</ID>
<type>DE_TO</type>
<position>177.5,-256.5</position>
<input>
<ID>IN_0</ID>735 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>1041</ID>
<type>DE_TO</type>
<position>177.5,-258.5</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>1042</ID>
<type>DE_TO</type>
<position>177.5,-260.5</position>
<input>
<ID>IN_0</ID>734 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>29.5,-238</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1043</ID>
<type>DE_TO</type>
<position>177.5,-262.5</position>
<input>
<ID>IN_0</ID>724 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>29.5,-241.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1044</ID>
<type>DE_TO</type>
<position>177.5,-248.5</position>
<input>
<ID>IN_0</ID>740 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>1045</ID>
<type>DE_TO</type>
<position>177.5,-250.5</position>
<input>
<ID>IN_0</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_LABEL</type>
<position>33,-192.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1046</ID>
<type>DE_TO</type>
<position>177.5,-252.5</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_LABEL</type>
<position>33,-196</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1047</ID>
<type>DE_TO</type>
<position>177.5,-254.5</position>
<input>
<ID>IN_0</ID>736 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_LABEL</type>
<position>33,-199.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1048</ID>
<type>AA_LABEL</type>
<position>115.5,-229</position>
<gparam>LABEL_TEXT Dez</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>270</ID>
<type>AA_LABEL</type>
<position>33,-203</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1049</ID>
<type>AA_LABEL</type>
<position>117,-248</position>
<gparam>LABEL_TEXT Unidade</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>AA_LABEL</type>
<position>33,-206.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>272</ID>
<type>AA_LABEL</type>
<position>33,-210</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1051</ID>
<type>AE_REGISTER8</type>
<position>167,-256</position>
<input>
<ID>IN_0</ID>730 </input>
<input>
<ID>IN_1</ID>731 </input>
<input>
<ID>IN_2</ID>732 </input>
<input>
<ID>IN_3</ID>737 </input>
<input>
<ID>IN_4</ID>741 </input>
<input>
<ID>IN_5</ID>742 </input>
<input>
<ID>IN_6</ID>743 </input>
<input>
<ID>IN_7</ID>744 </input>
<output>
<ID>OUT_0</ID>724 </output>
<output>
<ID>OUT_1</ID>734 </output>
<output>
<ID>OUT_2</ID>733 </output>
<output>
<ID>OUT_3</ID>735 </output>
<output>
<ID>OUT_4</ID>736 </output>
<output>
<ID>OUT_5</ID>738 </output>
<output>
<ID>OUT_6</ID>739 </output>
<output>
<ID>OUT_7</ID>740 </output>
<input>
<ID>clock</ID>746 </input>
<input>
<ID>load</ID>745 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_LABEL</type>
<position>33,-213.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>274</ID>
<type>AA_LABEL</type>
<position>33,-217</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>275</ID>
<type>AA_LABEL</type>
<position>33,-220.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>276</ID>
<type>AA_LABEL</type>
<position>33,-224</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>277</ID>
<type>AA_LABEL</type>
<position>33,-227.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>667</ID>
<type>AA_AND2</type>
<position>315,-269.5</position>
<input>
<ID>IN_0</ID>583 </input>
<input>
<ID>IN_1</ID>584 </input>
<output>
<ID>OUT</ID>585 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_LABEL</type>
<position>33,-231</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>668</ID>
<type>DA_FROM</type>
<position>307,-267.5</position>
<input>
<ID>IN_0</ID>583 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g0</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_LABEL</type>
<position>33,-234.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>669</ID>
<type>DA_FROM</type>
<position>307,-271.5</position>
<input>
<ID>IN_0</ID>584 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_LABEL</type>
<position>33,-238</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>670</ID>
<type>GA_LED</type>
<position>318.5,-283.5</position>
<input>
<ID>N_in0</ID>585 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>281</ID>
<type>AA_LABEL</type>
<position>33,-241.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>288</ID>
<type>AA_LABEL</type>
<position>59,-172.5</position>
<gparam>LABEL_TEXT G = X AND Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>GA_LED</type>
<position>48,-178</position>
<input>
<ID>N_in0</ID>320 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>290</ID>
<type>BI_DECODER_4x16</type>
<position>24.5,-173.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>231 </input>
<input>
<ID>IN_2</ID>230 </input>
<input>
<ID>IN_3</ID>265 </input>
<output>
<ID>OUT_0</ID>286 </output>
<output>
<ID>OUT_1</ID>314 </output>
<output>
<ID>OUT_10</ID>326 </output>
<output>
<ID>OUT_11</ID>325 </output>
<output>
<ID>OUT_12</ID>142 </output>
<output>
<ID>OUT_13</ID>143 </output>
<output>
<ID>OUT_14</ID>144 </output>
<output>
<ID>OUT_15</ID>145 </output>
<output>
<ID>OUT_2</ID>316 </output>
<output>
<ID>OUT_3</ID>317 </output>
<output>
<ID>OUT_4</ID>318 </output>
<output>
<ID>OUT_5</ID>319 </output>
<output>
<ID>OUT_6</ID>320 </output>
<output>
<ID>OUT_7</ID>321 </output>
<output>
<ID>OUT_8</ID>322 </output>
<output>
<ID>OUT_9</ID>324 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>291</ID>
<type>AA_LABEL</type>
<position>57.5,-155.5</position>
<gparam>LABEL_TEXT G = NOT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>AA_LABEL</type>
<position>58.5,-170</position>
<gparam>LABEL_TEXT G = X OR Y </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_LABEL</type>
<position>59,-167.5</position>
<gparam>LABEL_TEXT G = X XOR Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_LABEL</type>
<position>60,-164.5</position>
<gparam>LABEL_TEXT G = X XNOR Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>AA_LABEL</type>
<position>59,-158.5</position>
<gparam>LABEL_TEXT G = X NOR Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>297</ID>
<type>GA_LED</type>
<position>48,-175.5</position>
<input>
<ID>N_in0</ID>321 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>299</ID>
<type>GA_LED</type>
<position>48,-173</position>
<input>
<ID>N_in0</ID>322 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>301</ID>
<type>GA_LED</type>
<position>48,-190.5</position>
<input>
<ID>N_in0</ID>314 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>303</ID>
<type>GA_LED</type>
<position>48,-170.5</position>
<input>
<ID>N_in0</ID>324 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>316</ID>
<type>GA_LED</type>
<position>48,-168</position>
<input>
<ID>N_in0</ID>326 </input>
<input>
<ID>N_in3</ID>326 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>328</ID>
<type>GA_LED</type>
<position>48,-165</position>
<input>
<ID>N_in0</ID>325 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>329</ID>
<type>DA_FROM</type>
<position>13.5,-182.5</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>348</ID>
<type>AA_LABEL</type>
<position>60,-161.5</position>
<gparam>LABEL_TEXT G = X NAND Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>349</ID>
<type>GA_LED</type>
<position>48,-188</position>
<input>
<ID>N_in0</ID>316 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>DA_FROM</type>
<position>13.5,-177.5</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>351</ID>
<type>DA_FROM</type>
<position>13.5,-180</position>
<input>
<ID>IN_0</ID>231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>362</ID>
<type>DA_FROM</type>
<position>13.5,-175</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>363</ID>
<type>GA_LED</type>
<position>48,-185.5</position>
<input>
<ID>N_in0</ID>317 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>162.5,-196.5</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<wire>
<ID>772</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,-283.5,235,-283.5</points>
<connection>
<GID>1207</GID>
<name>N_in0</name></connection>
<intersection>235 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>235,-283.5,235,-269.5</points>
<connection>
<GID>1204</GID>
<name>OUT</name></connection>
<intersection>-283.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>773</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>210,-268.5,212.5,-268.5</points>
<connection>
<GID>1322</GID>
<name>IN_0</name></connection>
<intersection>210 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>210,-268.5,210,-267.5</points>
<intersection>-268.5 1</intersection>
<intersection>-267.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>209.5,-267.5,210,-267.5</points>
<connection>
<GID>1323</GID>
<name>IN_0</name></connection>
<intersection>210 5</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-190.5,137.5,-173.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_0</name></connection>
<intersection>-190.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>121,-190.5,137.5,-190.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-188.5,136.5,-172.5</points>
<intersection>-188.5 2</intersection>
<intersection>-172.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,-172.5,137.5,-172.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_1</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-188.5,136.5,-188.5</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>775</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-271.5,210,-270.5</points>
<intersection>-271.5 4</intersection>
<intersection>-270.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>210,-270.5,212.5,-270.5</points>
<connection>
<GID>1322</GID>
<name>IN_1</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>209.5,-271.5,210,-271.5</points>
<connection>
<GID>1324</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-186.5,135.5,-171.5</points>
<intersection>-186.5 2</intersection>
<intersection>-171.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-171.5,137.5,-171.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_2</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-186.5,135.5,-186.5</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>309.5,-268.5,312,-268.5</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>309.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>309.5,-268.5,309.5,-267.5</points>
<intersection>-268.5 1</intersection>
<intersection>-267.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>309,-267.5,309.5,-267.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>309.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-184.5,134.5,-170.5</points>
<intersection>-184.5 2</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134.5,-170.5,137.5,-170.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_3</name></connection>
<intersection>134.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-184.5,134.5,-184.5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>134.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,-271.5,309.5,-270.5</points>
<intersection>-271.5 4</intersection>
<intersection>-270.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>309.5,-270.5,312,-270.5</points>
<connection>
<GID>667</GID>
<name>IN_1</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>309,-271.5,309.5,-271.5</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118.5,-169.5,137.5,-169.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_4</name></connection>
<intersection>118.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>118.5,-171,118.5,-169.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-169.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>317.5,-283.5,318,-283.5</points>
<connection>
<GID>670</GID>
<name>N_in0</name></connection>
<intersection>318 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>318,-283.5,318,-269.5</points>
<connection>
<GID>667</GID>
<name>OUT</name></connection>
<intersection>-283.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118.5,-168.5,137.5,-168.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_5</name></connection>
<intersection>118.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>118.5,-169,118.5,-168.5</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>-168.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118.5,-167.5,137.5,-167.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_6</name></connection>
<intersection>118.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>118.5,-167.5,118.5,-167</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>-167.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-193.5,170.5,-190</points>
<intersection>-193.5 4</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>169.5,-190,170.5,-190</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>170.5,-193.5,174,-193.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>176,-144,192.5,-144</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>192.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192.5,-145,192.5,-144</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-144 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>184,-155,217.5,-155</points>
<intersection>184 5</intersection>
<intersection>192.5 4</intersection>
<intersection>217.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>217.5,-155,217.5,-153</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-155 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>192.5,-155,192.5,-148</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>-155 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>184,-155,184,-148</points>
<connection>
<GID>11</GID>
<name>CLK</name></connection>
<intersection>-155 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,-148,201.5,-146.5</points>
<intersection>-148 2</intersection>
<intersection>-146.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201.5,-146.5,205,-146.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198.5,-148,201.5,-148</points>
<connection>
<GID>6</GID>
<name>OUTINV_0</name></connection>
<intersection>201.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>211,-145.5,213,-145.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>213 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>213,-145.5,213,-145</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-145.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-145,198.5,-142.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-142.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198.5,-142.5,199.5,-142.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204,-144.5,204,-142.5</points>
<intersection>-144.5 1</intersection>
<intersection>-142.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204,-144.5,205,-144.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>204 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-142.5,204,-142.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>204 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118.5,-166.5,137.5,-166.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_7</name></connection>
<intersection>118.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>118.5,-166.5,118.5,-165</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>-166.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-165.5,134,-153.5</points>
<intersection>-165.5 1</intersection>
<intersection>-153.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-165.5,137.5,-165.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_8</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-153.5,134,-153.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-164.5,135,-151.5</points>
<intersection>-164.5 1</intersection>
<intersection>-151.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-164.5,137.5,-164.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_9</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-151.5,135,-151.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-163.5,136,-149.5</points>
<intersection>-163.5 1</intersection>
<intersection>-149.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-163.5,137.5,-163.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_10</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-149.5,136,-149.5</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-162.5,137,-147.5</points>
<intersection>-162.5 1</intersection>
<intersection>-147.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-162.5,137.5,-162.5</points>
<connection>
<GID>5</GID>
<name>ADDRESS_11</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-147.5,137,-147.5</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-190,154,-179</points>
<connection>
<GID>5</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-190 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-190,161.5,-190</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>154 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-189,153,-179</points>
<connection>
<GID>5</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-189 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153,-189,161.5,-189</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>153 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-188,152,-179</points>
<connection>
<GID>5</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-188 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152,-188,161.5,-188</points>
<connection>
<GID>137</GID>
<name>IN_2</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,-189.5,172.5,-188</points>
<intersection>-189.5 1</intersection>
<intersection>-188 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,-189.5,174,-189.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>172.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>169.5,-188,172.5,-188</points>
<connection>
<GID>137</GID>
<name>OUT_2</name></connection>
<intersection>172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,-191.5,171.5,-189</points>
<intersection>-191.5 2</intersection>
<intersection>-189 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-189,171.5,-189</points>
<connection>
<GID>137</GID>
<name>OUT_1</name></connection>
<intersection>171.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171.5,-191.5,174,-191.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173.5,-187.5,174,-187.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>173.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>173.5,-187.5,173.5,-187</points>
<intersection>-187.5 1</intersection>
<intersection>-187 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>169.5,-187,173.5,-187</points>
<connection>
<GID>137</GID>
<name>OUT_3</name></connection>
<intersection>173.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>169.5,-186,173.5,-186</points>
<connection>
<GID>137</GID>
<name>OUT_4</name></connection>
<intersection>173.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>173.5,-186,173.5,-185.5</points>
<intersection>-186 2</intersection>
<intersection>-185.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>173.5,-185.5,174,-185.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>173.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-187,151,-179</points>
<connection>
<GID>5</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-187 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-187,161.5,-187</points>
<connection>
<GID>137</GID>
<name>IN_3</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,-185,172.5,-183.5</points>
<intersection>-185 1</intersection>
<intersection>-183.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-185,172.5,-185</points>
<connection>
<GID>137</GID>
<name>OUT_5</name></connection>
<intersection>172.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172.5,-183.5,174,-183.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,-184,171.5,-181.5</points>
<intersection>-184 2</intersection>
<intersection>-181.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171.5,-181.5,174,-181.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>171.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169.5,-184,171.5,-184</points>
<connection>
<GID>137</GID>
<name>OUT_6</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-183,170.5,-179.5</points>
<intersection>-183 1</intersection>
<intersection>-179.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-183,170.5,-183</points>
<connection>
<GID>137</GID>
<name>OUT_7</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170.5,-179.5,174,-179.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-179,21.5,-179</points>
<connection>
<GID>290</GID>
<name>IN_2</name></connection>
<intersection>16.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>16.5,-179,16.5,-177.5</points>
<intersection>-179 1</intersection>
<intersection>-177.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>15.5,-177.5,16.5,-177.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>16.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-180,21.5,-180</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<connection>
<GID>351</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>810</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-283.5,218.5,-283.5</points>
<connection>
<GID>1325</GID>
<name>N_in0</name></connection>
<intersection>218.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>218.5,-283.5,218.5,-269.5</points>
<connection>
<GID>1322</GID>
<name>OUT</name></connection>
<intersection>-283.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-186,150,-179</points>
<connection>
<GID>5</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-186,161.5,-186</points>
<connection>
<GID>137</GID>
<name>IN_4</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>811</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>193.5,-268.5,196,-268.5</points>
<connection>
<GID>1214</GID>
<name>IN_0</name></connection>
<intersection>193.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>193.5,-268.5,193.5,-267.5</points>
<intersection>-268.5 1</intersection>
<intersection>-267.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>193,-267.5,193.5,-267.5</points>
<connection>
<GID>1309</GID>
<name>IN_0</name></connection>
<intersection>193.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>812</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,-271.5,193.5,-270.5</points>
<intersection>-271.5 4</intersection>
<intersection>-270.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>193.5,-270.5,196,-270.5</points>
<connection>
<GID>1214</GID>
<name>IN_1</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>193,-271.5,193.5,-271.5</points>
<connection>
<GID>1319</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>813</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>201.5,-283.5,202,-283.5</points>
<connection>
<GID>1320</GID>
<name>N_in0</name></connection>
<intersection>202 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>202,-283.5,202,-269.5</points>
<connection>
<GID>1214</GID>
<name>OUT</name></connection>
<intersection>-283.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-185,149,-179</points>
<connection>
<GID>5</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149,-185,161.5,-185</points>
<connection>
<GID>137</GID>
<name>IN_5</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-184,148,-179</points>
<connection>
<GID>5</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-184 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148,-184,161.5,-184</points>
<connection>
<GID>137</GID>
<name>IN_6</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,-183,147,-179</points>
<connection>
<GID>5</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-183 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-183,161.5,-183</points>
<connection>
<GID>137</GID>
<name>IN_7</name></connection>
<intersection>147 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>8</ID>
<points>17,-178,17,-175</points>
<intersection>-178 12</intersection>
<intersection>-175 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>17,-178,21.5,-178</points>
<connection>
<GID>290</GID>
<name>IN_3</name></connection>
<intersection>17 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>15.5,-175,17,-175</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>17 8</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>94.5,-203.5,95,-203.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>95 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>95,-203.5,95,-203.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-203.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-203.5,80.5,-203.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>65.5,-203.5,66,-203.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>66 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>66,-203.5,66,-203.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-203.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-193,39,-181</points>
<intersection>-193 1</intersection>
<intersection>-181 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-193,47,-193</points>
<connection>
<GID>250</GID>
<name>N_in0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-181,39,-181</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-181,164.5,-178</points>
<connection>
<GID>137</GID>
<name>load</name></connection>
<intersection>-178 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164,-178,164.5,-178</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-222,60,-222</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<connection>
<GID>531</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-229,60,-229</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<connection>
<GID>813</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-241.5,60,-241.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<connection>
<GID>815</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-259.5,139,-242.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_0</name></connection>
<intersection>-259.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-259.5,139,-259.5</points>
<connection>
<GID>1035</GID>
<name>OUT_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-235.5,60,-235.5</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<connection>
<GID>607</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-257.5,138,-241.5</points>
<intersection>-257.5 2</intersection>
<intersection>-241.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-241.5,139,-241.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_1</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-257.5,138,-257.5</points>
<connection>
<GID>1035</GID>
<name>OUT_1</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-196.5,164.5,-192</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<connection>
<GID>137</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-240.5,227,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_11</name></connection>
<intersection>-240.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,-240.5,230.5,-240.5</points>
<connection>
<GID>429</GID>
<name>IN_3</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-241.5,228,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_10</name></connection>
<intersection>-241.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228,-241.5,230.5,-241.5</points>
<connection>
<GID>429</GID>
<name>IN_2</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-242.5,229,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_9</name></connection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,-242.5,230.5,-242.5</points>
<connection>
<GID>429</GID>
<name>IN_1</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-243.5,230,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_8</name></connection>
<intersection>-243.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>230,-243.5,230.5,-243.5</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-182.5,17,-181</points>
<intersection>-182.5 8</intersection>
<intersection>-181 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>17,-181,21.5,-181</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>15.5,-182.5,17,-182.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-190.5,40,-180</points>
<intersection>-190.5 1</intersection>
<intersection>-180 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-190.5,47,-190.5</points>
<connection>
<GID>301</GID>
<name>N_in0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27.5,-180,40,-180</points>
<connection>
<GID>290</GID>
<name>OUT_1</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-188,47,-188</points>
<connection>
<GID>349</GID>
<name>N_in0</name></connection>
<intersection>41 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41,-188,41,-179</points>
<intersection>-188 1</intersection>
<intersection>-179 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>27.5,-179,41,-179</points>
<connection>
<GID>290</GID>
<name>OUT_2</name></connection>
<intersection>41 3</intersection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-185.5,42,-178</points>
<intersection>-185.5 1</intersection>
<intersection>-178 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-185.5,47,-185.5</points>
<connection>
<GID>363</GID>
<name>N_in0</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-178,42,-178</points>
<connection>
<GID>290</GID>
<name>OUT_3</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-183,47,-183</points>
<connection>
<GID>253</GID>
<name>N_in0</name></connection>
<intersection>43 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>43,-183,43,-177</points>
<intersection>-183 1</intersection>
<intersection>-177 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>27.5,-177,43,-177</points>
<connection>
<GID>290</GID>
<name>OUT_4</name></connection>
<intersection>43 5</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>27.5,-176.5,44,-176.5</points>
<intersection>27.5 8</intersection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-180.5,44,-176.5</points>
<intersection>-180.5 9</intersection>
<intersection>-176.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>27.5,-176.5,27.5,-176</points>
<connection>
<GID>290</GID>
<name>OUT_5</name></connection>
<intersection>-176.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>44,-180.5,47,-180.5</points>
<connection>
<GID>255</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-178,47,-178</points>
<connection>
<GID>289</GID>
<name>N_in0</name></connection>
<intersection>45 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>45,-178,45,-175</points>
<intersection>-178 1</intersection>
<intersection>-175 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>27.5,-175,45,-175</points>
<connection>
<GID>290</GID>
<name>OUT_6</name></connection>
<intersection>45 13</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-175.5,45.5,-174</points>
<intersection>-175.5 1</intersection>
<intersection>-174 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-175.5,47,-175.5</points>
<connection>
<GID>297</GID>
<name>N_in0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-174,45.5,-174</points>
<connection>
<GID>290</GID>
<name>OUT_7</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-173,47,-173</points>
<connection>
<GID>299</GID>
<name>N_in0</name></connection>
<connection>
<GID>290</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-172,44.5,-170.5</points>
<intersection>-172 2</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-170.5,47,-170.5</points>
<connection>
<GID>303</GID>
<name>N_in0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-172,44.5,-172</points>
<connection>
<GID>290</GID>
<name>OUT_9</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-170,43.5,-165</points>
<intersection>-170 2</intersection>
<intersection>-165 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-170,43.5,-170</points>
<connection>
<GID>290</GID>
<name>OUT_11</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-165,47,-165</points>
<connection>
<GID>328</GID>
<name>N_in0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-168,48,-168</points>
<connection>
<GID>316</GID>
<name>N_in0</name></connection>
<intersection>44 6</intersection>
<intersection>48 9</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>44,-171,44,-168</points>
<intersection>-171 8</intersection>
<intersection>-168 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>27.5,-171,44,-171</points>
<connection>
<GID>290</GID>
<name>OUT_10</name></connection>
<intersection>44 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>48,-168,48,-167</points>
<connection>
<GID>316</GID>
<name>N_in3</name></connection>
<intersection>-168 1</intersection></vsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-255.5,137,-240.5</points>
<intersection>-255.5 2</intersection>
<intersection>-240.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-240.5,139,-240.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_2</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-255.5,137,-255.5</points>
<connection>
<GID>1035</GID>
<name>OUT_2</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-253.5,136,-239.5</points>
<intersection>-253.5 2</intersection>
<intersection>-239.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-239.5,139,-239.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_3</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-253.5,136,-253.5</points>
<connection>
<GID>1035</GID>
<name>OUT_3</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-238.5,139,-238.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_4</name></connection>
<intersection>120 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>120,-240,120,-238.5</points>
<connection>
<GID>1034</GID>
<name>OUT_0</name></connection>
<intersection>-238.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-169,42.5,-162</points>
<intersection>-169 2</intersection>
<intersection>-162 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-162,47,-162</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-169,42.5,-169</points>
<connection>
<GID>290</GID>
<name>OUT_12</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-237.5,139,-237.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_5</name></connection>
<intersection>120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>120,-238,120,-237.5</points>
<connection>
<GID>1034</GID>
<name>OUT_1</name></connection>
<intersection>-237.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-168,41,-159</points>
<intersection>-168 2</intersection>
<intersection>-159 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-159,47,-159</points>
<connection>
<GID>151</GID>
<name>N_in0</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-168,41,-168</points>
<connection>
<GID>290</GID>
<name>OUT_13</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-236.5,139,-236.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_6</name></connection>
<intersection>120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>120,-236.5,120,-236</points>
<connection>
<GID>1034</GID>
<name>OUT_2</name></connection>
<intersection>-236.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-167,40,-156</points>
<intersection>-167 2</intersection>
<intersection>-156 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-156,47,-156</points>
<connection>
<GID>152</GID>
<name>N_in0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-167,40,-167</points>
<connection>
<GID>290</GID>
<name>OUT_14</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-262.5,172,-259</points>
<intersection>-262.5 4</intersection>
<intersection>-259 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>171,-259,172,-259</points>
<connection>
<GID>1051</GID>
<name>OUT_0</name></connection>
<intersection>172 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>172,-262.5,175.5,-262.5</points>
<connection>
<GID>1043</GID>
<name>IN_0</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-166,38.5,-153</points>
<intersection>-166 2</intersection>
<intersection>-153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-153,47,-153</points>
<connection>
<GID>153</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-166,38.5,-166</points>
<connection>
<GID>290</GID>
<name>OUT_15</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231,-237.5,231,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-237.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>231,-237.5,247.5,-237.5</points>
<connection>
<GID>428</GID>
<name>IN_7</name></connection>
<intersection>231 0</intersection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-235.5,139,-235.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_7</name></connection>
<intersection>120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>120,-235.5,120,-234</points>
<connection>
<GID>1034</GID>
<name>OUT_3</name></connection>
<intersection>-235.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-236.5,232,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-236.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232,-236.5,245.5,-236.5</points>
<intersection>232 0</intersection>
<intersection>245.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>245.5,-238.5,245.5,-236.5</points>
<intersection>-238.5 6</intersection>
<intersection>-236.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>245.5,-238.5,247.5,-238.5</points>
<connection>
<GID>428</GID>
<name>IN_6</name></connection>
<intersection>245.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-234.5,135.5,-222.5</points>
<intersection>-234.5 1</intersection>
<intersection>-222.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-234.5,139,-234.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_8</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-222.5,135.5,-222.5</points>
<connection>
<GID>1037</GID>
<name>OUT_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-235.5,233,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233,-235.5,244.5,-235.5</points>
<intersection>233 0</intersection>
<intersection>244.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>244.5,-239.5,244.5,-235.5</points>
<intersection>-239.5 5</intersection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>244.5,-239.5,247.5,-239.5</points>
<connection>
<GID>428</GID>
<name>IN_5</name></connection>
<intersection>244.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-233.5,136.5,-220.5</points>
<intersection>-233.5 1</intersection>
<intersection>-220.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,-233.5,139,-233.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_9</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-220.5,136.5,-220.5</points>
<connection>
<GID>1037</GID>
<name>OUT_1</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,-234.5,234,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-234.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,-234.5,243.5,-234.5</points>
<intersection>234 0</intersection>
<intersection>243.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>243.5,-240.5,243.5,-234.5</points>
<intersection>-240.5 6</intersection>
<intersection>-234.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>243.5,-240.5,247.5,-240.5</points>
<connection>
<GID>428</GID>
<name>IN_4</name></connection>
<intersection>243.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-232.5,137.5,-218.5</points>
<intersection>-232.5 1</intersection>
<intersection>-218.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,-232.5,139,-232.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_10</name></connection>
<intersection>137.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-218.5,137.5,-218.5</points>
<connection>
<GID>1037</GID>
<name>OUT_2</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,-233.5,235,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-233.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,-233.5,242.5,-233.5</points>
<intersection>235 0</intersection>
<intersection>242.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>242.5,-241.5,242.5,-233.5</points>
<intersection>-241.5 6</intersection>
<intersection>-233.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>242.5,-241.5,247.5,-241.5</points>
<connection>
<GID>428</GID>
<name>IN_3</name></connection>
<intersection>242.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-231.5,138.5,-216.5</points>
<intersection>-231.5 1</intersection>
<intersection>-216.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-231.5,139,-231.5</points>
<connection>
<GID>1036</GID>
<name>ADDRESS_11</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-216.5,138.5,-216.5</points>
<connection>
<GID>1037</GID>
<name>OUT_3</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-232.5,236,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-232.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,-232.5,241.5,-232.5</points>
<intersection>236 0</intersection>
<intersection>241.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>241.5,-242.5,241.5,-232.5</points>
<intersection>-242.5 6</intersection>
<intersection>-232.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>241.5,-242.5,247.5,-242.5</points>
<connection>
<GID>428</GID>
<name>IN_2</name></connection>
<intersection>241.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-259,155.5,-248</points>
<connection>
<GID>1036</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-259 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,-259,163,-259</points>
<connection>
<GID>1051</GID>
<name>IN_0</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-231.5,237,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-231.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>237,-231.5,240.5,-231.5</points>
<intersection>237 0</intersection>
<intersection>240.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>240.5,-243.5,240.5,-231.5</points>
<intersection>-243.5 6</intersection>
<intersection>-231.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>240.5,-243.5,247.5,-243.5</points>
<connection>
<GID>428</GID>
<name>IN_1</name></connection>
<intersection>240.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-258,154.5,-248</points>
<connection>
<GID>1036</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-258 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154.5,-258,163,-258</points>
<connection>
<GID>1051</GID>
<name>IN_1</name></connection>
<intersection>154.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-230.5,238,-229</points>
<connection>
<GID>160</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-230.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238,-230.5,239.5,-230.5</points>
<intersection>238 0</intersection>
<intersection>239.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>239.5,-244.5,239.5,-230.5</points>
<intersection>-244.5 6</intersection>
<intersection>-230.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>239.5,-244.5,247.5,-244.5</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>239.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-257,153.5,-248</points>
<connection>
<GID>1036</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-257 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153.5,-257,163,-257</points>
<connection>
<GID>1051</GID>
<name>IN_2</name></connection>
<intersection>153.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-258.5,174,-257</points>
<intersection>-258.5 1</intersection>
<intersection>-257 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,-258.5,175.5,-258.5</points>
<connection>
<GID>1041</GID>
<name>IN_0</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>171,-257,174,-257</points>
<connection>
<GID>1051</GID>
<name>OUT_2</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-227,208,-223.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>-227 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>198,-227,208,-227</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-260.5,173,-258</points>
<intersection>-260.5 2</intersection>
<intersection>-258 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-258,173,-258</points>
<connection>
<GID>1051</GID>
<name>OUT_1</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>173,-260.5,175.5,-260.5</points>
<connection>
<GID>1042</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206,-225,206,-222.5</points>
<intersection>-225 2</intersection>
<intersection>-222.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206,-222.5,208,-222.5</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>206 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198,-225,206,-225</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>206 0</intersection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>175,-256.5,175.5,-256.5</points>
<connection>
<GID>1040</GID>
<name>IN_0</name></connection>
<intersection>175 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>175,-256.5,175,-256</points>
<intersection>-256.5 1</intersection>
<intersection>-256 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>171,-256,175,-256</points>
<connection>
<GID>1051</GID>
<name>OUT_3</name></connection>
<intersection>175 12</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-221.5,208,-221.5</points>
<connection>
<GID>169</GID>
<name>IN_2</name></connection>
<intersection>198 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>198,-223,198,-221.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-221.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>171,-255,175,-255</points>
<connection>
<GID>1051</GID>
<name>OUT_4</name></connection>
<intersection>175 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>175,-255,175,-254.5</points>
<intersection>-255 2</intersection>
<intersection>-254.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>175,-254.5,175.5,-254.5</points>
<connection>
<GID>1047</GID>
<name>IN_0</name></connection>
<intersection>175 5</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>12</ID>
<points>198,-221,198,-220.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-220.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>198,-220.5,208,-220.5</points>
<connection>
<GID>169</GID>
<name>IN_3</name></connection>
<intersection>198 12</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-256,152.5,-248</points>
<connection>
<GID>1036</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-256 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152.5,-256,163,-256</points>
<connection>
<GID>1051</GID>
<name>IN_3</name></connection>
<intersection>152.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-219.5,208,-219.5</points>
<connection>
<GID>169</GID>
<name>IN_4</name></connection>
<intersection>198 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>198,-219.5,198,-219</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>-219.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-254,174,-252.5</points>
<intersection>-254 1</intersection>
<intersection>-252.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-254,174,-254</points>
<connection>
<GID>1051</GID>
<name>OUT_5</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,-252.5,175.5,-252.5</points>
<connection>
<GID>1046</GID>
<name>IN_0</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-218.5,208,-218.5</points>
<connection>
<GID>169</GID>
<name>IN_5</name></connection>
<intersection>198 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>198,-218.5,198,-217</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-218.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-253,173,-250.5</points>
<intersection>-253 2</intersection>
<intersection>-250.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173,-250.5,175.5,-250.5</points>
<connection>
<GID>1045</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171,-253,173,-253</points>
<connection>
<GID>1051</GID>
<name>OUT_6</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206,-217.5,206,-215</points>
<intersection>-217.5 1</intersection>
<intersection>-215 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206,-217.5,208,-217.5</points>
<connection>
<GID>169</GID>
<name>IN_6</name></connection>
<intersection>206 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198,-215,206,-215</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>206 0</intersection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-252,172,-248.5</points>
<intersection>-252 1</intersection>
<intersection>-248.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-252,172,-252</points>
<connection>
<GID>1051</GID>
<name>OUT_7</name></connection>
<intersection>172 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-248.5,175.5,-248.5</points>
<connection>
<GID>1044</GID>
<name>IN_0</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-213,208,-213</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>208 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>208,-216.5,208,-213</points>
<connection>
<GID>169</GID>
<name>IN_7</name></connection>
<intersection>-213 1</intersection></vsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-255,151.5,-248</points>
<connection>
<GID>1036</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-255 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,-255,163,-255</points>
<connection>
<GID>1051</GID>
<name>IN_4</name></connection>
<intersection>151.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211,-230,211,-225.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<connection>
<GID>169</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-254,150.5,-248</points>
<connection>
<GID>1036</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-254 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-254,163,-254</points>
<connection>
<GID>1051</GID>
<name>IN_5</name></connection>
<intersection>150.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>211,-214.5,211,-212.5</points>
<connection>
<GID>169</GID>
<name>load</name></connection>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-253,149.5,-248</points>
<connection>
<GID>1036</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-253 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-253,163,-253</points>
<connection>
<GID>1051</GID>
<name>IN_6</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-223.5,221.5,-223.5</points>
<connection>
<GID>160</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-252,148.5,-248</points>
<connection>
<GID>1036</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-252 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148.5,-252,163,-252</points>
<connection>
<GID>1051</GID>
<name>IN_7</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-222.5,221.5,-222.5</points>
<connection>
<GID>160</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>169</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-221.5,221.5,-221.5</points>
<connection>
<GID>160</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>169</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-250,166,-247</points>
<connection>
<GID>1051</GID>
<name>load</name></connection>
<intersection>-247 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165.5,-247,166,-247</points>
<connection>
<GID>1181</GID>
<name>IN_0</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-220.5,221.5,-220.5</points>
<connection>
<GID>160</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>169</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-265.5,166,-261</points>
<connection>
<GID>1182</GID>
<name>IN_0</name></connection>
<connection>
<GID>1051</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>51,-203.5,51.5,-203.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<connection>
<GID>227</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-219.5,221.5,-219.5</points>
<connection>
<GID>160</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>169</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>293,-268.5,295.5,-268.5</points>
<connection>
<GID>1189</GID>
<name>IN_0</name></connection>
<intersection>293 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>293,-268.5,293,-267.5</points>
<intersection>-268.5 1</intersection>
<intersection>-267.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>292.5,-267.5,293,-267.5</points>
<connection>
<GID>1190</GID>
<name>IN_0</name></connection>
<intersection>293 5</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-218.5,221.5,-218.5</points>
<connection>
<GID>160</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>169</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-217.5,221.5,-217.5</points>
<connection>
<GID>160</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>169</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-216.5,221.5,-216.5</points>
<connection>
<GID>160</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>169</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>758</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-271.5,293,-270.5</points>
<intersection>-271.5 4</intersection>
<intersection>-270.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-270.5,295.5,-270.5</points>
<connection>
<GID>1189</GID>
<name>IN_1</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>292.5,-271.5,293,-271.5</points>
<connection>
<GID>1191</GID>
<name>IN_0</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>301,-283.5,301.5,-283.5</points>
<connection>
<GID>1192</GID>
<name>N_in0</name></connection>
<intersection>301.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>301.5,-283.5,301.5,-269.5</points>
<connection>
<GID>1189</GID>
<name>OUT</name></connection>
<intersection>-283.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,-268.5,279,-268.5</points>
<connection>
<GID>1199</GID>
<name>IN_0</name></connection>
<intersection>276.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>276.5,-268.5,276.5,-267.5</points>
<intersection>-268.5 1</intersection>
<intersection>-267.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>276,-267.5,276.5,-267.5</points>
<connection>
<GID>1200</GID>
<name>IN_0</name></connection>
<intersection>276.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276.5,-271.5,276.5,-270.5</points>
<intersection>-271.5 4</intersection>
<intersection>-270.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>276.5,-270.5,279,-270.5</points>
<connection>
<GID>1199</GID>
<name>IN_1</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>276,-271.5,276.5,-271.5</points>
<connection>
<GID>1201</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>284.5,-283.5,285,-283.5</points>
<connection>
<GID>1202</GID>
<name>N_in0</name></connection>
<intersection>285 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>285,-283.5,285,-269.5</points>
<connection>
<GID>1199</GID>
<name>OUT</name></connection>
<intersection>-283.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>260,-268.5,262.5,-268.5</points>
<connection>
<GID>1194</GID>
<name>IN_0</name></connection>
<intersection>260 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>260,-268.5,260,-267.5</points>
<intersection>-268.5 1</intersection>
<intersection>-267.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>259.5,-267.5,260,-267.5</points>
<connection>
<GID>1195</GID>
<name>IN_0</name></connection>
<intersection>260 5</intersection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-271.5,260,-270.5</points>
<intersection>-271.5 4</intersection>
<intersection>-270.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>260,-270.5,262.5,-270.5</points>
<connection>
<GID>1194</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>259.5,-271.5,260,-271.5</points>
<connection>
<GID>1196</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>268,-283.5,268.5,-283.5</points>
<connection>
<GID>1197</GID>
<name>N_in0</name></connection>
<intersection>268.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>268.5,-283.5,268.5,-269.5</points>
<connection>
<GID>1194</GID>
<name>OUT</name></connection>
<intersection>-283.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243,-268.5,245.5,-268.5</points>
<connection>
<GID>1209</GID>
<name>IN_0</name></connection>
<intersection>243 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>243,-268.5,243,-267.5</points>
<intersection>-268.5 1</intersection>
<intersection>-267.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>242.5,-267.5,243,-267.5</points>
<connection>
<GID>1210</GID>
<name>IN_0</name></connection>
<intersection>243 5</intersection></hsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-271.5,243,-270.5</points>
<intersection>-271.5 4</intersection>
<intersection>-270.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>243,-270.5,245.5,-270.5</points>
<connection>
<GID>1209</GID>
<name>IN_1</name></connection>
<intersection>243 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>242.5,-271.5,243,-271.5</points>
<connection>
<GID>1211</GID>
<name>IN_0</name></connection>
<intersection>243 0</intersection></hsegment></shape></wire>
<wire>
<ID>769</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>251,-283.5,251.5,-283.5</points>
<connection>
<GID>1212</GID>
<name>N_in0</name></connection>
<intersection>251.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>251.5,-283.5,251.5,-269.5</points>
<connection>
<GID>1209</GID>
<name>OUT</name></connection>
<intersection>-283.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>770</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>226.5,-268.5,229,-268.5</points>
<connection>
<GID>1204</GID>
<name>IN_0</name></connection>
<intersection>226.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>226.5,-268.5,226.5,-267.5</points>
<intersection>-268.5 1</intersection>
<intersection>-267.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>226,-267.5,226.5,-267.5</points>
<connection>
<GID>1205</GID>
<name>IN_0</name></connection>
<intersection>226.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>771</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-271.5,226.5,-270.5</points>
<intersection>-271.5 4</intersection>
<intersection>-270.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-270.5,229,-270.5</points>
<connection>
<GID>1204</GID>
<name>IN_1</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226,-271.5,226.5,-271.5</points>
<connection>
<GID>1206</GID>
<name>IN_0</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>491.528,2408.83,722.497,2290.75</PageViewport>
<gate>
<ID>595</ID>
<type>AA_AND3</type>
<position>708.5,2378</position>
<input>
<ID>IN_0</ID>699 </input>
<input>
<ID>IN_1</ID>700 </input>
<input>
<ID>IN_2</ID>701 </input>
<output>
<ID>OUT</ID>697 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>596</ID>
<type>AA_LABEL</type>
<position>685.5,2389</position>
<gparam>LABEL_TEXT Complemento de 2 de Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>597</ID>
<type>AI_INVERTER_4BIT</type>
<position>669,2378</position>
<input>
<ID>IN_0</ID>612 </input>
<input>
<ID>IN_1</ID>613 </input>
<input>
<ID>IN_2</ID>614 </input>
<input>
<ID>IN_3</ID>615 </input>
<output>
<ID>OUT_0</ID>622 </output>
<output>
<ID>OUT_1</ID>623 </output>
<output>
<ID>OUT_2</ID>624 </output>
<output>
<ID>OUT_3</ID>625 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>598</ID>
<type>AI_INVERTER_4BIT</type>
<position>669,2373.5</position>
<input>
<ID>IN_0</ID>608 </input>
<input>
<ID>IN_1</ID>609 </input>
<input>
<ID>IN_2</ID>610 </input>
<input>
<ID>IN_3</ID>611 </input>
<output>
<ID>OUT_0</ID>618 </output>
<output>
<ID>OUT_1</ID>619 </output>
<output>
<ID>OUT_2</ID>620 </output>
<output>
<ID>OUT_3</ID>621 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>599</ID>
<type>DA_FROM</type>
<position>659,2377</position>
<input>
<ID>IN_0</ID>612 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>603</ID>
<type>DA_FROM</type>
<position>659,2374.5</position>
<input>
<ID>IN_0</ID>611 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>605</ID>
<type>DA_FROM</type>
<position>659,2372</position>
<input>
<ID>IN_0</ID>610 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>609</ID>
<type>DA_FROM</type>
<position>659,2369.5</position>
<input>
<ID>IN_0</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>610</ID>
<type>DA_FROM</type>
<position>659,2367</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>611</ID>
<type>DA_FROM</type>
<position>659,2384.5</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>612</ID>
<type>DA_FROM</type>
<position>659,2382</position>
<input>
<ID>IN_0</ID>614 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>613</ID>
<type>DA_FROM</type>
<position>659,2379.5</position>
<input>
<ID>IN_0</ID>613 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>816</ID>
<type>DE_TO</type>
<position>644,2323</position>
<input>
<ID>IN_0</ID>716 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as4</lparam></gate>
<gate>
<ID>624</ID>
<type>DE_TO</type>
<position>614.5,2332</position>
<input>
<ID>IN_0</ID>937 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cs</lparam></gate>
<gate>
<ID>625</ID>
<type>AE_FULLADDER_4BIT</type>
<position>680,2366.5</position>
<input>
<ID>IN_0</ID>621 </input>
<input>
<ID>IN_1</ID>620 </input>
<input>
<ID>IN_2</ID>619 </input>
<input>
<ID>IN_3</ID>618 </input>
<output>
<ID>OUT_0</ID>644 </output>
<output>
<ID>OUT_1</ID>645 </output>
<output>
<ID>OUT_2</ID>646 </output>
<output>
<ID>OUT_3</ID>647 </output>
<input>
<ID>carry_in</ID>616 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>818</ID>
<type>DE_TO</type>
<position>644,2320.5</position>
<input>
<ID>IN_0</ID>717 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as5</lparam></gate>
<gate>
<ID>626</ID>
<type>AE_FULLADDER_4BIT</type>
<position>698,2366.5</position>
<input>
<ID>IN_0</ID>625 </input>
<input>
<ID>IN_1</ID>624 </input>
<input>
<ID>IN_2</ID>623 </input>
<input>
<ID>IN_3</ID>622 </input>
<output>
<ID>OUT_0</ID>640 </output>
<output>
<ID>OUT_1</ID>641 </output>
<output>
<ID>OUT_2</ID>642 </output>
<output>
<ID>OUT_3</ID>643 </output>
<input>
<ID>carry_in</ID>935 </input>
<output>
<ID>carry_out</ID>616 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>627</ID>
<type>DE_TO</type>
<position>507,2354</position>
<input>
<ID>IN_0</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cix</lparam></gate>
<gate>
<ID>820</ID>
<type>DE_TO</type>
<position>644,2318</position>
<input>
<ID>IN_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as6</lparam></gate>
<gate>
<ID>628</ID>
<type>DE_TO</type>
<position>509,2308</position>
<input>
<ID>IN_0</ID>939 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cdx</lparam></gate>
<gate>
<ID>821</ID>
<type>DE_TO</type>
<position>644,2315.5</position>
<input>
<ID>IN_0</ID>749 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as7</lparam></gate>
<gate>
<ID>629</ID>
<type>DE_TO</type>
<position>561.5,2307.5</position>
<input>
<ID>IN_0</ID>940 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cdy</lparam></gate>
<gate>
<ID>1016</ID>
<type>AA_LABEL</type>
<position>598.5,2406</position>
<gparam>LABEL_TEXT Unidade Aritmetica</gparam>
<gparam>TEXT_HEIGHT 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>839</ID>
<type>DE_TO</type>
<position>644,2333</position>
<input>
<ID>IN_0</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as0</lparam></gate>
<gate>
<ID>840</ID>
<type>DE_TO</type>
<position>644,2330.5</position>
<input>
<ID>IN_0</ID>713 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as1</lparam></gate>
<gate>
<ID>842</ID>
<type>DE_TO</type>
<position>644,2328</position>
<input>
<ID>IN_0</ID>714 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as2</lparam></gate>
<gate>
<ID>843</ID>
<type>DE_TO</type>
<position>644,2325.5</position>
<input>
<ID>IN_0</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as3</lparam></gate>
<gate>
<ID>846</ID>
<type>EE_VDD</type>
<position>543,2366</position>
<output>
<ID>OUT_0</ID>933 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>847</ID>
<type>AE_FULLADDER_4BIT</type>
<position>516.5,2314.5</position>
<input>
<ID>IN_0</ID>757 </input>
<input>
<ID>IN_1</ID>759 </input>
<input>
<ID>IN_2</ID>750 </input>
<input>
<ID>IN_3</ID>751 </input>
<input>
<ID>IN_B_0</ID>884 </input>
<input>
<ID>IN_B_1</ID>884 </input>
<input>
<ID>IN_B_2</ID>884 </input>
<input>
<ID>IN_B_3</ID>884 </input>
<output>
<ID>OUT_0</ID>914 </output>
<output>
<ID>OUT_1</ID>915 </output>
<output>
<ID>OUT_2</ID>916 </output>
<output>
<ID>OUT_3</ID>917 </output>
<input>
<ID>carry_in</ID>752 </input>
<output>
<ID>carry_out</ID>939 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>848</ID>
<type>AE_FULLADDER_4BIT</type>
<position>534.5,2314.5</position>
<input>
<ID>IN_0</ID>753 </input>
<input>
<ID>IN_1</ID>754 </input>
<input>
<ID>IN_2</ID>755 </input>
<input>
<ID>IN_3</ID>756 </input>
<input>
<ID>IN_B_0</ID>884 </input>
<input>
<ID>IN_B_1</ID>884 </input>
<input>
<ID>IN_B_2</ID>884 </input>
<input>
<ID>IN_B_3</ID>884 </input>
<output>
<ID>OUT_0</ID>910 </output>
<output>
<ID>OUT_1</ID>911 </output>
<output>
<ID>OUT_2</ID>912 </output>
<output>
<ID>OUT_3</ID>913 </output>
<output>
<ID>carry_out</ID>752 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>849</ID>
<type>DA_FROM</type>
<position>509,2329.5</position>
<input>
<ID>IN_0</ID>756 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>850</ID>
<type>DA_FROM</type>
<position>509,2327</position>
<input>
<ID>IN_0</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>851</ID>
<type>DA_FROM</type>
<position>509,2324.5</position>
<input>
<ID>IN_0</ID>759 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>852</ID>
<type>DA_FROM</type>
<position>509,2322</position>
<input>
<ID>IN_0</ID>750 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>853</ID>
<type>DA_FROM</type>
<position>509,2319.5</position>
<input>
<ID>IN_0</ID>751 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>854</ID>
<type>DA_FROM</type>
<position>509,2337</position>
<input>
<ID>IN_0</ID>753 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>855</ID>
<type>DA_FROM</type>
<position>509,2334.5</position>
<input>
<ID>IN_0</ID>754 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>856</ID>
<type>DA_FROM</type>
<position>509,2332</position>
<input>
<ID>IN_0</ID>755 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>857</ID>
<type>EE_VDD</type>
<position>596.5,2369</position>
<output>
<ID>OUT_0</ID>934 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>859</ID>
<type>AE_FULLADDER_4BIT</type>
<position>570.5,2315.5</position>
<input>
<ID>IN_0</ID>821 </input>
<input>
<ID>IN_1</ID>822 </input>
<input>
<ID>IN_2</ID>814 </input>
<input>
<ID>IN_3</ID>815 </input>
<input>
<ID>IN_B_0</ID>851 </input>
<input>
<ID>IN_B_1</ID>851 </input>
<input>
<ID>IN_B_2</ID>851 </input>
<input>
<ID>IN_B_3</ID>851 </input>
<output>
<ID>OUT_0</ID>897 </output>
<output>
<ID>OUT_1</ID>898 </output>
<output>
<ID>OUT_2</ID>899 </output>
<output>
<ID>OUT_3</ID>900 </output>
<input>
<ID>carry_in</ID>816 </input>
<output>
<ID>carry_out</ID>940 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>860</ID>
<type>AE_FULLADDER_4BIT</type>
<position>588.5,2315.5</position>
<input>
<ID>IN_0</ID>817 </input>
<input>
<ID>IN_1</ID>818 </input>
<input>
<ID>IN_2</ID>819 </input>
<input>
<ID>IN_3</ID>820 </input>
<input>
<ID>IN_B_0</ID>851 </input>
<input>
<ID>IN_B_1</ID>851 </input>
<input>
<ID>IN_B_2</ID>851 </input>
<input>
<ID>IN_B_3</ID>851 </input>
<output>
<ID>OUT_0</ID>893 </output>
<output>
<ID>OUT_1</ID>894 </output>
<output>
<ID>OUT_2</ID>895 </output>
<output>
<ID>OUT_3</ID>896 </output>
<output>
<ID>carry_out</ID>816 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>861</ID>
<type>DA_FROM</type>
<position>563.5,2330.5</position>
<input>
<ID>IN_0</ID>820 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>862</ID>
<type>DA_FROM</type>
<position>563.5,2328</position>
<input>
<ID>IN_0</ID>821 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>863</ID>
<type>DA_FROM</type>
<position>563.5,2325.5</position>
<input>
<ID>IN_0</ID>822 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>671</ID>
<type>DE_TO</type>
<position>562,2354.5</position>
<input>
<ID>IN_0</ID>941 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ciy</lparam></gate>
<gate>
<ID>864</ID>
<type>DA_FROM</type>
<position>563.5,2323</position>
<input>
<ID>IN_0</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>865</ID>
<type>DA_FROM</type>
<position>563.5,2320.5</position>
<input>
<ID>IN_0</ID>815 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>673</ID>
<type>EE_VDD</type>
<position>707.5,2371.5</position>
<output>
<ID>OUT_0</ID>935 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>866</ID>
<type>DA_FROM</type>
<position>563.5,2338</position>
<input>
<ID>IN_0</ID>817 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>867</ID>
<type>DA_FROM</type>
<position>563.5,2335.5</position>
<input>
<ID>IN_0</ID>818 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>675</ID>
<type>AA_MUX_2x1</type>
<position>707.5,2360</position>
<input>
<ID>IN_0</ID>632 </input>
<input>
<ID>IN_1</ID>640 </input>
<output>
<ID>OUT</ID>649 </output>
<input>
<ID>SEL_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>868</ID>
<type>DA_FROM</type>
<position>563.5,2333</position>
<input>
<ID>IN_0</ID>819 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>676</ID>
<type>AA_LABEL</type>
<position>629,2389.5</position>
<gparam>LABEL_TEXT Adicao e Subtracao</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>869</ID>
<type>EE_VDD</type>
<position>539.5,2323</position>
<output>
<ID>OUT_0</ID>884 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>677</ID>
<type>DA_FROM</type>
<position>703,2380</position>
<input>
<ID>IN_0</ID>699 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>870</ID>
<type>EE_VDD</type>
<position>593.5,2325</position>
<output>
<ID>OUT_0</ID>851 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>678</ID>
<type>DA_FROM</type>
<position>703,2378</position>
<input>
<ID>IN_0</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>871</ID>
<type>DE_TO</type>
<position>592,2350.5</position>
<input>
<ID>IN_0</ID>889 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy3</lparam></gate>
<gate>
<ID>679</ID>
<type>AE_FULLADDER_4BIT</type>
<position>516,2362.5</position>
<input>
<ID>IN_0</ID>589 </input>
<input>
<ID>IN_1</ID>590 </input>
<input>
<ID>IN_2</ID>505 </input>
<input>
<ID>IN_3</ID>506 </input>
<output>
<ID>OUT_0</ID>905 </output>
<output>
<ID>OUT_1</ID>906 </output>
<output>
<ID>OUT_2</ID>909 </output>
<output>
<ID>OUT_3</ID>908 </output>
<input>
<ID>carry_in</ID>507 </input>
<output>
<ID>carry_out</ID>938 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>872</ID>
<type>DE_TO</type>
<position>592,2353</position>
<input>
<ID>IN_0</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy2</lparam></gate>
<gate>
<ID>680</ID>
<type>AE_FULLADDER_4BIT</type>
<position>534,2362.5</position>
<input>
<ID>IN_0</ID>512 </input>
<input>
<ID>IN_1</ID>586 </input>
<input>
<ID>IN_2</ID>587 </input>
<input>
<ID>IN_3</ID>588 </input>
<output>
<ID>OUT_0</ID>901 </output>
<output>
<ID>OUT_1</ID>902 </output>
<output>
<ID>OUT_2</ID>903 </output>
<output>
<ID>OUT_3</ID>904 </output>
<input>
<ID>carry_in</ID>933 </input>
<output>
<ID>carry_out</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>873</ID>
<type>DE_TO</type>
<position>592,2355.5</position>
<input>
<ID>IN_0</ID>891 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy1</lparam></gate>
<gate>
<ID>681</ID>
<type>AE_FULLADDER_4BIT</type>
<position>570,2363</position>
<input>
<ID>IN_0</ID>595 </input>
<input>
<ID>IN_1</ID>594 </input>
<input>
<ID>IN_2</ID>511 </input>
<input>
<ID>IN_3</ID>510 </input>
<output>
<ID>OUT_0</ID>888 </output>
<output>
<ID>OUT_1</ID>887 </output>
<output>
<ID>OUT_2</ID>886 </output>
<output>
<ID>OUT_3</ID>885 </output>
<input>
<ID>carry_in</ID>509 </input>
<output>
<ID>carry_out</ID>941 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>874</ID>
<type>DE_TO</type>
<position>592,2358</position>
<input>
<ID>IN_0</ID>892 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy0</lparam></gate>
<gate>
<ID>682</ID>
<type>AE_FULLADDER_4BIT</type>
<position>588,2363</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>598 </input>
<input>
<ID>IN_2</ID>597 </input>
<input>
<ID>IN_3</ID>596 </input>
<output>
<ID>OUT_0</ID>892 </output>
<output>
<ID>OUT_1</ID>891 </output>
<output>
<ID>OUT_2</ID>890 </output>
<output>
<ID>OUT_3</ID>889 </output>
<input>
<ID>carry_in</ID>934 </input>
<output>
<ID>carry_out</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>875</ID>
<type>DE_TO</type>
<position>592,2340.5</position>
<input>
<ID>IN_0</ID>885 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy7</lparam></gate>
<gate>
<ID>683</ID>
<type>DA_FROM</type>
<position>703,2376</position>
<input>
<ID>IN_0</ID>701 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>876</ID>
<type>DE_TO</type>
<position>592,2343</position>
<input>
<ID>IN_0</ID>886 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy6</lparam></gate>
<gate>
<ID>684</ID>
<type>AA_LABEL</type>
<position>521,2389.5</position>
<gparam>LABEL_TEXT Incremento e Decremento de X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>877</ID>
<type>DE_TO</type>
<position>592,2345.5</position>
<input>
<ID>IN_0</ID>887 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy5</lparam></gate>
<gate>
<ID>685</ID>
<type>AA_LABEL</type>
<position>576,2389.5</position>
<gparam>LABEL_TEXT Incremento e Decremento de Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>878</ID>
<type>DE_TO</type>
<position>592,2348</position>
<input>
<ID>IN_0</ID>888 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy4</lparam></gate>
<gate>
<ID>686</ID>
<type>AA_MUX_2x1</type>
<position>707.5,2355</position>
<input>
<ID>IN_0</ID>639 </input>
<input>
<ID>IN_1</ID>641 </input>
<output>
<ID>OUT</ID>651 </output>
<input>
<ID>SEL_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>879</ID>
<type>FF_GND</type>
<position>649.5,2336.5</position>
<output>
<ID>OUT_0</ID>932 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>687</ID>
<type>AA_MUX_2x1</type>
<position>707.5,2350</position>
<input>
<ID>IN_0</ID>638 </input>
<input>
<ID>IN_1</ID>642 </input>
<output>
<ID>OUT</ID>653 </output>
<input>
<ID>SEL_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>880</ID>
<type>DE_TO</type>
<position>592.5,2303</position>
<input>
<ID>IN_0</ID>896 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy3</lparam></gate>
<gate>
<ID>688</ID>
<type>AA_MUX_2x1</type>
<position>707.5,2345</position>
<input>
<ID>IN_0</ID>637 </input>
<input>
<ID>IN_1</ID>643 </input>
<output>
<ID>OUT</ID>670 </output>
<input>
<ID>SEL_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>689</ID>
<type>AA_MUX_2x1</type>
<position>707.5,2335</position>
<input>
<ID>IN_0</ID>635 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>652 </output>
<input>
<ID>SEL_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>690</ID>
<type>AA_MUX_2x1</type>
<position>707.5,2330</position>
<input>
<ID>IN_0</ID>634 </input>
<input>
<ID>IN_1</ID>646 </input>
<output>
<ID>OUT</ID>650 </output>
<input>
<ID>SEL_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>691</ID>
<type>AA_MUX_2x1</type>
<position>707.5,2325</position>
<input>
<ID>IN_0</ID>633 </input>
<input>
<ID>IN_1</ID>647 </input>
<output>
<ID>OUT</ID>648 </output>
<input>
<ID>SEL_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>692</ID>
<type>AA_MUX_2x1</type>
<position>707.5,2340</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>644 </input>
<output>
<ID>OUT</ID>659 </output>
<input>
<ID>SEL_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>885</ID>
<type>DE_TO</type>
<position>592.5,2305.5</position>
<input>
<ID>IN_0</ID>895 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy2</lparam></gate>
<gate>
<ID>693</ID>
<type>DA_FROM</type>
<position>702.5,2344</position>
<input>
<ID>IN_0</ID>637 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>886</ID>
<type>DE_TO</type>
<position>592.5,2308</position>
<input>
<ID>IN_0</ID>894 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy1</lparam></gate>
<gate>
<ID>694</ID>
<type>DA_FROM</type>
<position>702.5,2339</position>
<input>
<ID>IN_0</ID>636 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>887</ID>
<type>DE_TO</type>
<position>592.5,2310.5</position>
<input>
<ID>IN_0</ID>893 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy0</lparam></gate>
<gate>
<ID>695</ID>
<type>DA_FROM</type>
<position>702.5,2334</position>
<input>
<ID>IN_0</ID>635 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>888</ID>
<type>DE_TO</type>
<position>592.5,2293</position>
<input>
<ID>IN_0</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy7</lparam></gate>
<gate>
<ID>696</ID>
<type>DA_FROM</type>
<position>703,2329</position>
<input>
<ID>IN_0</ID>634 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>889</ID>
<type>DE_TO</type>
<position>592.5,2295.5</position>
<input>
<ID>IN_0</ID>899 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy6</lparam></gate>
<gate>
<ID>697</ID>
<type>DA_FROM</type>
<position>703,2324</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>890</ID>
<type>DE_TO</type>
<position>592.5,2298</position>
<input>
<ID>IN_0</ID>898 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy5</lparam></gate>
<gate>
<ID>891</ID>
<type>DE_TO</type>
<position>592.5,2300.5</position>
<input>
<ID>IN_0</ID>897 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy4</lparam></gate>
<gate>
<ID>892</ID>
<type>DE_TO</type>
<position>538,2350</position>
<input>
<ID>IN_0</ID>904 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx3</lparam></gate>
<gate>
<ID>700</ID>
<type>DA_FROM</type>
<position>702.5,2359</position>
<input>
<ID>IN_0</ID>632 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>893</ID>
<type>DE_TO</type>
<position>538,2352.5</position>
<input>
<ID>IN_0</ID>903 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx2</lparam></gate>
<gate>
<ID>894</ID>
<type>DE_TO</type>
<position>538,2355</position>
<input>
<ID>IN_0</ID>902 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx1</lparam></gate>
<gate>
<ID>895</ID>
<type>DE_TO</type>
<position>538,2357.5</position>
<input>
<ID>IN_0</ID>901 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx0</lparam></gate>
<gate>
<ID>896</ID>
<type>DE_TO</type>
<position>538,2340</position>
<input>
<ID>IN_0</ID>908 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx7</lparam></gate>
<gate>
<ID>897</ID>
<type>DE_TO</type>
<position>538,2342.5</position>
<input>
<ID>IN_0</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx6</lparam></gate>
<gate>
<ID>898</ID>
<type>DE_TO</type>
<position>538,2345</position>
<input>
<ID>IN_0</ID>906 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx5</lparam></gate>
<gate>
<ID>899</ID>
<type>DE_TO</type>
<position>538,2347.5</position>
<input>
<ID>IN_0</ID>905 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx4</lparam></gate>
<gate>
<ID>900</ID>
<type>DE_TO</type>
<position>538,2302</position>
<input>
<ID>IN_0</ID>913 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx3</lparam></gate>
<gate>
<ID>901</ID>
<type>DE_TO</type>
<position>538,2304.5</position>
<input>
<ID>IN_0</ID>912 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx2</lparam></gate>
<gate>
<ID>902</ID>
<type>DE_TO</type>
<position>538,2307</position>
<input>
<ID>IN_0</ID>911 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx1</lparam></gate>
<gate>
<ID>903</ID>
<type>DE_TO</type>
<position>538,2309.5</position>
<input>
<ID>IN_0</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx0</lparam></gate>
<gate>
<ID>904</ID>
<type>DE_TO</type>
<position>538,2292</position>
<input>
<ID>IN_0</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx7</lparam></gate>
<gate>
<ID>905</ID>
<type>DE_TO</type>
<position>538,2294.5</position>
<input>
<ID>IN_0</ID>916 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx6</lparam></gate>
<gate>
<ID>906</ID>
<type>DE_TO</type>
<position>538,2297</position>
<input>
<ID>IN_0</ID>915 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx5</lparam></gate>
<gate>
<ID>907</ID>
<type>DE_TO</type>
<position>538,2299.5</position>
<input>
<ID>IN_0</ID>914 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx4</lparam></gate>
<gate>
<ID>716</ID>
<type>DA_FROM</type>
<position>702.5,2354</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>717</ID>
<type>DA_FROM</type>
<position>702.5,2349</position>
<input>
<ID>IN_0</ID>638 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>719</ID>
<type>DA_FROM</type>
<position>508.5,2377.5</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>720</ID>
<type>DA_FROM</type>
<position>508.5,2375</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>721</ID>
<type>DE_TO</type>
<position>712.5,2345</position>
<input>
<ID>IN_0</ID>670 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'3</lparam></gate>
<gate>
<ID>722</ID>
<type>DA_FROM</type>
<position>508.5,2372.5</position>
<input>
<ID>IN_0</ID>590 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>723</ID>
<type>DE_TO</type>
<position>712.5,2350</position>
<input>
<ID>IN_0</ID>653 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'2</lparam></gate>
<gate>
<ID>543</ID>
<type>DA_FROM</type>
<position>562.5,2378</position>
<input>
<ID>IN_0</ID>596 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>740</ID>
<type>DA_FROM</type>
<position>508.5,2370</position>
<input>
<ID>IN_0</ID>505 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>741</ID>
<type>DE_TO</type>
<position>712.5,2355</position>
<input>
<ID>IN_0</ID>651 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'1</lparam></gate>
<gate>
<ID>548</ID>
<type>DA_FROM</type>
<position>562.5,2375.5</position>
<input>
<ID>IN_0</ID>595 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>742</ID>
<type>DA_FROM</type>
<position>508.5,2367.5</position>
<input>
<ID>IN_0</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>549</ID>
<type>DA_FROM</type>
<position>562.5,2373</position>
<input>
<ID>IN_0</ID>594 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>743</ID>
<type>DE_TO</type>
<position>712.5,2360</position>
<input>
<ID>IN_0</ID>649 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'0</lparam></gate>
<gate>
<ID>744</ID>
<type>DA_FROM</type>
<position>508.5,2385</position>
<input>
<ID>IN_0</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>745</ID>
<type>DE_TO</type>
<position>712.5,2325</position>
<input>
<ID>IN_0</ID>648 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'7</lparam></gate>
<gate>
<ID>746</ID>
<type>DA_FROM</type>
<position>508.5,2382.5</position>
<input>
<ID>IN_0</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>553</ID>
<type>DA_FROM</type>
<position>562.5,2370.5</position>
<input>
<ID>IN_0</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>747</ID>
<type>DE_TO</type>
<position>712.5,2330</position>
<input>
<ID>IN_0</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'6</lparam></gate>
<gate>
<ID>748</ID>
<type>DA_FROM</type>
<position>508.5,2380</position>
<input>
<ID>IN_0</ID>587 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>749</ID>
<type>DE_TO</type>
<position>712.5,2335</position>
<input>
<ID>IN_0</ID>652 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'5</lparam></gate>
<gate>
<ID>750</ID>
<type>DE_TO</type>
<position>712.5,2340</position>
<input>
<ID>IN_0</ID>659 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'4</lparam></gate>
<gate>
<ID>751</ID>
<type>AE_FULLADDER_4BIT</type>
<position>622,2338</position>
<input>
<ID>IN_0</ID>692 </input>
<input>
<ID>IN_1</ID>693 </input>
<input>
<ID>IN_2</ID>671 </input>
<input>
<ID>IN_3</ID>672 </input>
<input>
<ID>IN_B_0</ID>617 </input>
<input>
<ID>IN_B_1</ID>593 </input>
<input>
<ID>IN_B_2</ID>592 </input>
<input>
<ID>IN_B_3</ID>591 </input>
<output>
<ID>OUT_0</ID>716 </output>
<output>
<ID>OUT_1</ID>717 </output>
<output>
<ID>OUT_2</ID>718 </output>
<output>
<ID>OUT_3</ID>749 </output>
<input>
<ID>carry_in</ID>673 </input>
<output>
<ID>carry_out</ID>937 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>752</ID>
<type>AE_FULLADDER_4BIT</type>
<position>640,2338</position>
<input>
<ID>IN_0</ID>674 </input>
<input>
<ID>IN_1</ID>675 </input>
<input>
<ID>IN_2</ID>676 </input>
<input>
<ID>IN_3</ID>691 </input>
<input>
<ID>IN_B_0</ID>627 </input>
<input>
<ID>IN_B_1</ID>628 </input>
<input>
<ID>IN_B_2</ID>629 </input>
<input>
<ID>IN_B_3</ID>626 </input>
<output>
<ID>OUT_0</ID>712 </output>
<output>
<ID>OUT_1</ID>713 </output>
<output>
<ID>OUT_2</ID>714 </output>
<output>
<ID>OUT_3</ID>715 </output>
<input>
<ID>carry_in</ID>932 </input>
<output>
<ID>carry_out</ID>673 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>753</ID>
<type>DA_FROM</type>
<position>614.5,2354</position>
<input>
<ID>IN_0</ID>691 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>754</ID>
<type>DA_FROM</type>
<position>614.5,2351.5</position>
<input>
<ID>IN_0</ID>692 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>755</ID>
<type>DA_FROM</type>
<position>614.5,2349</position>
<input>
<ID>IN_0</ID>693 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>756</ID>
<type>DA_FROM</type>
<position>614.5,2346.5</position>
<input>
<ID>IN_0</ID>671 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>757</ID>
<type>DA_FROM</type>
<position>614.5,2344</position>
<input>
<ID>IN_0</ID>672 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>758</ID>
<type>DA_FROM</type>
<position>614.5,2361.5</position>
<input>
<ID>IN_0</ID>674 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>759</ID>
<type>DA_FROM</type>
<position>614.5,2359</position>
<input>
<ID>IN_0</ID>675 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>760</ID>
<type>DA_FROM</type>
<position>614.5,2356.5</position>
<input>
<ID>IN_0</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>761</ID>
<type>DA_FROM</type>
<position>614.5,2376</position>
<input>
<ID>IN_0</ID>626 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'3</lparam></gate>
<gate>
<ID>762</ID>
<type>DA_FROM</type>
<position>614.5,2373.5</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'4</lparam></gate>
<gate>
<ID>763</ID>
<type>DA_FROM</type>
<position>614.5,2371</position>
<input>
<ID>IN_0</ID>593 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'5</lparam></gate>
<gate>
<ID>764</ID>
<type>DA_FROM</type>
<position>614.5,2368.5</position>
<input>
<ID>IN_0</ID>592 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'6</lparam></gate>
<gate>
<ID>571</ID>
<type>DA_FROM</type>
<position>562.5,2368</position>
<input>
<ID>IN_0</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>765</ID>
<type>DA_FROM</type>
<position>614.5,2366</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'7</lparam></gate>
<gate>
<ID>572</ID>
<type>DA_FROM</type>
<position>562.5,2385.5</position>
<input>
<ID>IN_0</ID>599 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>766</ID>
<type>DA_FROM</type>
<position>614.5,2383.5</position>
<input>
<ID>IN_0</ID>627 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'0</lparam></gate>
<gate>
<ID>573</ID>
<type>DA_FROM</type>
<position>562.5,2383</position>
<input>
<ID>IN_0</ID>598 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>767</ID>
<type>DA_FROM</type>
<position>614.5,2381</position>
<input>
<ID>IN_0</ID>628 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'1</lparam></gate>
<gate>
<ID>768</ID>
<type>DA_FROM</type>
<position>614.5,2378.5</position>
<input>
<ID>IN_0</ID>629 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y'2</lparam></gate>
<gate>
<ID>575</ID>
<type>DA_FROM</type>
<position>562.5,2380.5</position>
<input>
<ID>IN_0</ID>597 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<wire>
<ID>586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>531,2366.5,531,2382.5</points>
<connection>
<GID>680</GID>
<name>IN_1</name></connection>
<intersection>2382.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,2382.5,531,2382.5</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>531 0</intersection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530,2366.5,530,2380</points>
<connection>
<GID>680</GID>
<name>IN_2</name></connection>
<intersection>2380 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,2380,530,2380</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>530 0</intersection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>529,2366.5,529,2377.5</points>
<connection>
<GID>680</GID>
<name>IN_3</name></connection>
<intersection>2377.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,2377.5,529,2377.5</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>529 0</intersection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,2366.5,514,2375</points>
<connection>
<GID>679</GID>
<name>IN_0</name></connection>
<intersection>2375 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,2375,514,2375</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513,2366.5,513,2372.5</points>
<connection>
<GID>679</GID>
<name>IN_1</name></connection>
<intersection>2372.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,2372.5,513,2372.5</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>513 0</intersection></hsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>624,2342,624,2366</points>
<connection>
<GID>751</GID>
<name>IN_B_3</name></connection>
<intersection>2366 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2366,624,2366</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>624 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>625,2342,625,2368.5</points>
<connection>
<GID>751</GID>
<name>IN_B_2</name></connection>
<intersection>2368.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2368.5,625,2368.5</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>625 0</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>626,2342,626,2371</points>
<connection>
<GID>751</GID>
<name>IN_B_1</name></connection>
<intersection>2371 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2371,626,2371</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>626 0</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>567,2367,567,2373</points>
<connection>
<GID>681</GID>
<name>IN_1</name></connection>
<intersection>2373 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>564.5,2373,567,2373</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>567 2</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>568,2367,568,2375.5</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<intersection>2375.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>564.5,2375.5,568,2375.5</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>568 0</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>564.5,2378,583,2378</points>
<connection>
<GID>543</GID>
<name>IN_0</name></connection>
<intersection>583 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>583,2367,583,2378</points>
<connection>
<GID>682</GID>
<name>IN_3</name></connection>
<intersection>2378 1</intersection></vsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584,2367,584,2380.5</points>
<connection>
<GID>682</GID>
<name>IN_2</name></connection>
<intersection>2380.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>564.5,2380.5,584,2380.5</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>584 0</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585,2367,585,2383</points>
<connection>
<GID>682</GID>
<name>IN_1</name></connection>
<intersection>2383 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>564.5,2383,585,2383</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>585 0</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>564.5,2385.5,586,2385.5</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>586 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>586,2367,586,2385.5</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>2385.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667,2367,667,2372</points>
<connection>
<GID>598</GID>
<name>IN_0</name></connection>
<intersection>2367 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>661,2367,667,2367</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<intersection>667 0</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666,2369.5,666,2373</points>
<intersection>2369.5 2</intersection>
<intersection>2373 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>666,2373,667,2373</points>
<connection>
<GID>598</GID>
<name>IN_1</name></connection>
<intersection>666 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>661,2369.5,666,2369.5</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<intersection>666 0</intersection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>665,2372,665,2374</points>
<intersection>2372 2</intersection>
<intersection>2374 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>665,2374,667,2374</points>
<connection>
<GID>598</GID>
<name>IN_2</name></connection>
<intersection>665 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>661,2372,665,2372</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>665 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,2374.5,667,2374.5</points>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>667 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>667,2374.5,667,2375</points>
<connection>
<GID>598</GID>
<name>IN_3</name></connection>
<intersection>2374.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,2377,667,2377</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>667 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>667,2376.5,667,2377</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>2377 1</intersection></vsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>665,2377.5,667,2377.5</points>
<connection>
<GID>597</GID>
<name>IN_1</name></connection>
<intersection>665 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>665,2377.5,665,2379.5</points>
<intersection>2377.5 1</intersection>
<intersection>2379.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>661,2379.5,665,2379.5</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>665 3</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666,2378.5,666,2382</points>
<intersection>2378.5 2</intersection>
<intersection>2382 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>661,2382,666,2382</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>666 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>666,2378.5,667,2378.5</points>
<connection>
<GID>597</GID>
<name>IN_2</name></connection>
<intersection>666 0</intersection></hsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667,2379.5,667,2384.5</points>
<connection>
<GID>597</GID>
<name>IN_3</name></connection>
<intersection>2384.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>661,2384.5,667,2384.5</points>
<connection>
<GID>611</GID>
<name>IN_0</name></connection>
<intersection>667 0</intersection></hsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,2367.5,690,2367.5</points>
<connection>
<GID>625</GID>
<name>carry_in</name></connection>
<connection>
<GID>626</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>627,2342,627,2373.5</points>
<connection>
<GID>751</GID>
<name>IN_B_0</name></connection>
<intersection>2373.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2373.5,627,2373.5</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>627 0</intersection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>675,2370.5,675,2372</points>
<connection>
<GID>625</GID>
<name>IN_3</name></connection>
<intersection>2372 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>671,2372,675,2372</points>
<connection>
<GID>598</GID>
<name>OUT_0</name></connection>
<intersection>675 0</intersection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>676,2370.5,676,2373</points>
<connection>
<GID>625</GID>
<name>IN_2</name></connection>
<intersection>2373 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>671,2373,676,2373</points>
<connection>
<GID>598</GID>
<name>OUT_1</name></connection>
<intersection>676 0</intersection></hsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>677,2370.5,677,2374</points>
<connection>
<GID>625</GID>
<name>IN_1</name></connection>
<intersection>2374 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>671,2374,677,2374</points>
<connection>
<GID>598</GID>
<name>OUT_2</name></connection>
<intersection>677 0</intersection></hsegment></shape></wire>
<wire>
<ID>814</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>566.5,2319.5,566.5,2323</points>
<connection>
<GID>859</GID>
<name>IN_2</name></connection>
<intersection>2323 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>565.5,2323,566.5,2323</points>
<connection>
<GID>864</GID>
<name>IN_0</name></connection>
<intersection>566.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>678,2370.5,678,2375</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>2375 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>671,2375,678,2375</points>
<connection>
<GID>598</GID>
<name>OUT_3</name></connection>
<intersection>678 0</intersection></hsegment></shape></wire>
<wire>
<ID>815</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>565.5,2319.5,565.5,2320.5</points>
<connection>
<GID>865</GID>
<name>IN_0</name></connection>
<connection>
<GID>859</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>693,2370.5,693,2376.5</points>
<connection>
<GID>626</GID>
<name>IN_3</name></connection>
<intersection>2376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>671,2376.5,693,2376.5</points>
<connection>
<GID>597</GID>
<name>OUT_0</name></connection>
<intersection>693 0</intersection></hsegment></shape></wire>
<wire>
<ID>816</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>578.5,2316.5,580.5,2316.5</points>
<connection>
<GID>859</GID>
<name>carry_in</name></connection>
<connection>
<GID>860</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>694,2370.5,694,2377.5</points>
<connection>
<GID>626</GID>
<name>IN_2</name></connection>
<intersection>2377.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>671,2377.5,694,2377.5</points>
<connection>
<GID>597</GID>
<name>OUT_1</name></connection>
<intersection>694 0</intersection></hsegment></shape></wire>
<wire>
<ID>817</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586.5,2319.5,586.5,2338</points>
<connection>
<GID>860</GID>
<name>IN_0</name></connection>
<intersection>2338 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>565.5,2338,586.5,2338</points>
<connection>
<GID>866</GID>
<name>IN_0</name></connection>
<intersection>586.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>695,2370.5,695,2378.5</points>
<connection>
<GID>626</GID>
<name>IN_1</name></connection>
<intersection>2378.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>671,2378.5,695,2378.5</points>
<connection>
<GID>597</GID>
<name>OUT_2</name></connection>
<intersection>695 0</intersection></hsegment></shape></wire>
<wire>
<ID>818</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,2319.5,585.5,2335.5</points>
<connection>
<GID>860</GID>
<name>IN_1</name></connection>
<intersection>2335.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>565.5,2335.5,585.5,2335.5</points>
<connection>
<GID>867</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>696,2370.5,696,2379.5</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>2379.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>671,2379.5,696,2379.5</points>
<connection>
<GID>597</GID>
<name>OUT_3</name></connection>
<intersection>696 0</intersection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>642,2342,642,2376</points>
<connection>
<GID>752</GID>
<name>IN_B_3</name></connection>
<intersection>2376 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2376,642,2376</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>642 0</intersection></hsegment></shape></wire>
<wire>
<ID>819</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584.5,2319.5,584.5,2333</points>
<connection>
<GID>860</GID>
<name>IN_2</name></connection>
<intersection>2333 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>565.5,2333,584.5,2333</points>
<connection>
<GID>868</GID>
<name>IN_0</name></connection>
<intersection>584.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>645,2342,645,2383.5</points>
<connection>
<GID>752</GID>
<name>IN_B_0</name></connection>
<intersection>2383.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2383.5,645,2383.5</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>645 0</intersection></hsegment></shape></wire>
<wire>
<ID>820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,2319.5,583.5,2330.5</points>
<connection>
<GID>860</GID>
<name>IN_3</name></connection>
<intersection>2330.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>565.5,2330.5,583.5,2330.5</points>
<connection>
<GID>861</GID>
<name>IN_0</name></connection>
<intersection>583.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644,2342,644,2381</points>
<connection>
<GID>752</GID>
<name>IN_B_1</name></connection>
<intersection>2381 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2381,644,2381</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<intersection>644 0</intersection></hsegment></shape></wire>
<wire>
<ID>821</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>568.5,2319.5,568.5,2328</points>
<connection>
<GID>859</GID>
<name>IN_0</name></connection>
<intersection>2328 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>565.5,2328,568.5,2328</points>
<connection>
<GID>862</GID>
<name>IN_0</name></connection>
<intersection>568.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>643,2342,643,2378.5</points>
<connection>
<GID>752</GID>
<name>IN_B_2</name></connection>
<intersection>2378.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2378.5,643,2378.5</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>643 0</intersection></hsegment></shape></wire>
<wire>
<ID>822</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>567.5,2319.5,567.5,2325.5</points>
<connection>
<GID>859</GID>
<name>IN_1</name></connection>
<intersection>2325.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>565.5,2325.5,567.5,2325.5</points>
<connection>
<GID>863</GID>
<name>IN_0</name></connection>
<intersection>567.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>704.5,2359,705.5,2359</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<connection>
<GID>700</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>705,2324,705.5,2324</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<connection>
<GID>697</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>705,2329,705.5,2329</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<connection>
<GID>696</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>704.5,2334,705.5,2334</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<connection>
<GID>695</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>704.5,2339,705.5,2339</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<connection>
<GID>694</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>704.5,2344,705.5,2344</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<connection>
<GID>693</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>704.5,2349,705.5,2349</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<connection>
<GID>717</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>704.5,2354,705.5,2354</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<connection>
<GID>716</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>699.5,2361,699.5,2362.5</points>
<connection>
<GID>626</GID>
<name>OUT_0</name></connection>
<intersection>2361 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>699.5,2361,705.5,2361</points>
<connection>
<GID>675</GID>
<name>IN_1</name></connection>
<intersection>699.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>698.5,2356,698.5,2362.5</points>
<connection>
<GID>626</GID>
<name>OUT_1</name></connection>
<intersection>2356 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>698.5,2356,705.5,2356</points>
<connection>
<GID>686</GID>
<name>IN_1</name></connection>
<intersection>698.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697.5,2351,697.5,2362.5</points>
<connection>
<GID>626</GID>
<name>OUT_2</name></connection>
<intersection>2351 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>697.5,2351,705.5,2351</points>
<connection>
<GID>687</GID>
<name>IN_1</name></connection>
<intersection>697.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>696.5,2346,696.5,2362.5</points>
<connection>
<GID>626</GID>
<name>OUT_3</name></connection>
<intersection>2346 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>696.5,2346,705.5,2346</points>
<connection>
<GID>688</GID>
<name>IN_1</name></connection>
<intersection>696.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>681.5,2341,681.5,2362.5</points>
<connection>
<GID>625</GID>
<name>OUT_0</name></connection>
<intersection>2341 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>681.5,2341,705.5,2341</points>
<connection>
<GID>692</GID>
<name>IN_1</name></connection>
<intersection>681.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,2336,680.5,2362.5</points>
<connection>
<GID>625</GID>
<name>OUT_1</name></connection>
<intersection>2336 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680.5,2336,705.5,2336</points>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>679.5,2331,679.5,2362.5</points>
<connection>
<GID>625</GID>
<name>OUT_2</name></connection>
<intersection>2331 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>679.5,2331,705.5,2331</points>
<connection>
<GID>690</GID>
<name>IN_1</name></connection>
<intersection>679.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>678.5,2326,678.5,2362.5</points>
<connection>
<GID>625</GID>
<name>OUT_3</name></connection>
<intersection>2326 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>678.5,2326,705.5,2326</points>
<connection>
<GID>691</GID>
<name>IN_1</name></connection>
<intersection>678.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>709.5,2325,710.5,2325</points>
<connection>
<GID>691</GID>
<name>OUT</name></connection>
<connection>
<GID>745</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>709.5,2360,710.5,2360</points>
<connection>
<GID>675</GID>
<name>OUT</name></connection>
<connection>
<GID>743</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>709.5,2330,710.5,2330</points>
<connection>
<GID>690</GID>
<name>OUT</name></connection>
<connection>
<GID>747</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>709.5,2355,710.5,2355</points>
<connection>
<GID>686</GID>
<name>OUT</name></connection>
<connection>
<GID>741</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>709.5,2335,710.5,2335</points>
<connection>
<GID>689</GID>
<name>OUT</name></connection>
<connection>
<GID>749</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>709.5,2350,710.5,2350</points>
<connection>
<GID>687</GID>
<name>OUT</name></connection>
<connection>
<GID>723</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>851</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593.5,2319.5,593.5,2324</points>
<connection>
<GID>870</GID>
<name>OUT_0</name></connection>
<connection>
<GID>860</GID>
<name>IN_B_0</name></connection>
<intersection>2322.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>572.5,2322.5,593.5,2322.5</points>
<intersection>572.5 7</intersection>
<intersection>573.5 12</intersection>
<intersection>574.5 14</intersection>
<intersection>575.5 11</intersection>
<intersection>590.5 16</intersection>
<intersection>591.5 20</intersection>
<intersection>592.5 8</intersection>
<intersection>593.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>572.5,2319.5,572.5,2322.5</points>
<connection>
<GID>859</GID>
<name>IN_B_3</name></connection>
<intersection>2322.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>592.5,2319.5,592.5,2322.5</points>
<connection>
<GID>860</GID>
<name>IN_B_1</name></connection>
<intersection>2322.5 5</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>575.5,2319.5,575.5,2322.5</points>
<connection>
<GID>859</GID>
<name>IN_B_0</name></connection>
<intersection>2322.5 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>573.5,2319.5,573.5,2322.5</points>
<connection>
<GID>859</GID>
<name>IN_B_2</name></connection>
<intersection>2322.5 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>574.5,2319.5,574.5,2322.5</points>
<connection>
<GID>859</GID>
<name>IN_B_1</name></connection>
<intersection>2322.5 5</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>590.5,2319.5,590.5,2322.5</points>
<connection>
<GID>860</GID>
<name>IN_B_3</name></connection>
<intersection>2322.5 5</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>591.5,2319.5,591.5,2322.5</points>
<connection>
<GID>860</GID>
<name>IN_B_2</name></connection>
<intersection>2322.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>709.5,2340,710.5,2340</points>
<connection>
<GID>692</GID>
<name>OUT</name></connection>
<connection>
<GID>750</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>709.5,2345,710.5,2345</points>
<connection>
<GID>688</GID>
<name>OUT</name></connection>
<connection>
<GID>721</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618,2342,618,2346.5</points>
<connection>
<GID>751</GID>
<name>IN_2</name></connection>
<intersection>2346.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2346.5,618,2346.5</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<intersection>618 0</intersection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>617,2342,617,2344</points>
<connection>
<GID>751</GID>
<name>IN_3</name></connection>
<intersection>2344 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>616.5,2344,617,2344</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>617 0</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>630,2339,632,2339</points>
<connection>
<GID>751</GID>
<name>carry_in</name></connection>
<connection>
<GID>752</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>638,2342,638,2361.5</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>2361.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2361.5,638,2361.5</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<intersection>638 0</intersection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>637,2342,637,2359</points>
<connection>
<GID>752</GID>
<name>IN_1</name></connection>
<intersection>2359 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2359,637,2359</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>637 0</intersection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>636,2342,636,2356.5</points>
<connection>
<GID>752</GID>
<name>IN_2</name></connection>
<intersection>2356.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2356.5,636,2356.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>636 0</intersection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>635,2342,635,2354</points>
<connection>
<GID>752</GID>
<name>IN_3</name></connection>
<intersection>2354 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2354,635,2354</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<intersection>635 0</intersection></hsegment></shape></wire>
<wire>
<ID>884</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539.5,2318.5,539.5,2322</points>
<connection>
<GID>869</GID>
<name>OUT_0</name></connection>
<connection>
<GID>848</GID>
<name>IN_B_0</name></connection>
<intersection>2321 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>518.5,2321,539.5,2321</points>
<intersection>518.5 10</intersection>
<intersection>519.5 11</intersection>
<intersection>520.5 12</intersection>
<intersection>521.5 13</intersection>
<intersection>536.5 14</intersection>
<intersection>537.5 15</intersection>
<intersection>538.5 16</intersection>
<intersection>539.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>518.5,2318.5,518.5,2321</points>
<connection>
<GID>847</GID>
<name>IN_B_3</name></connection>
<intersection>2321 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>519.5,2318.5,519.5,2321</points>
<connection>
<GID>847</GID>
<name>IN_B_2</name></connection>
<intersection>2321 2</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>520.5,2318.5,520.5,2321</points>
<connection>
<GID>847</GID>
<name>IN_B_1</name></connection>
<intersection>2321 2</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>521.5,2318.5,521.5,2321</points>
<connection>
<GID>847</GID>
<name>IN_B_0</name></connection>
<intersection>2321 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>536.5,2318.5,536.5,2321</points>
<connection>
<GID>848</GID>
<name>IN_B_3</name></connection>
<intersection>2321 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>537.5,2318.5,537.5,2321</points>
<connection>
<GID>848</GID>
<name>IN_B_2</name></connection>
<intersection>2321 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>538.5,2318.5,538.5,2321</points>
<connection>
<GID>848</GID>
<name>IN_B_1</name></connection>
<intersection>2321 2</intersection></vsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>620,2342,620,2351.5</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>2351.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>616.5,2351.5,620,2351.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>620 0</intersection></hsegment></shape></wire>
<wire>
<ID>885</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>568.5,2340.5,568.5,2359</points>
<connection>
<GID>681</GID>
<name>OUT_3</name></connection>
<intersection>2340.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>568.5,2340.5,590,2340.5</points>
<connection>
<GID>875</GID>
<name>IN_0</name></connection>
<intersection>568.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>619,2342,619,2349</points>
<connection>
<GID>751</GID>
<name>IN_1</name></connection>
<intersection>2349 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,2349,619,2349</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<intersection>619 0</intersection></hsegment></shape></wire>
<wire>
<ID>886</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>569.5,2343,569.5,2359</points>
<connection>
<GID>681</GID>
<name>OUT_2</name></connection>
<intersection>2343 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>569.5,2343,590,2343</points>
<connection>
<GID>876</GID>
<name>IN_0</name></connection>
<intersection>569.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>887</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>570.5,2345.5,570.5,2359</points>
<connection>
<GID>681</GID>
<name>OUT_1</name></connection>
<intersection>2345.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>570.5,2345.5,590,2345.5</points>
<connection>
<GID>877</GID>
<name>IN_0</name></connection>
<intersection>570.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>888</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,2348,571.5,2359</points>
<connection>
<GID>681</GID>
<name>OUT_0</name></connection>
<intersection>2348 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>571.5,2348,590,2348</points>
<connection>
<GID>878</GID>
<name>IN_0</name></connection>
<intersection>571.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>889</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586.5,2350.5,586.5,2359</points>
<connection>
<GID>682</GID>
<name>OUT_3</name></connection>
<intersection>2350.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>586.5,2350.5,590,2350.5</points>
<connection>
<GID>871</GID>
<name>IN_0</name></connection>
<intersection>586.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>890</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587.5,2353,587.5,2359</points>
<connection>
<GID>682</GID>
<name>OUT_2</name></connection>
<intersection>2353 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>587.5,2353,590,2353</points>
<connection>
<GID>872</GID>
<name>IN_0</name></connection>
<intersection>587.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>711.5,2378,716.5,2378</points>
<connection>
<GID>595</GID>
<name>OUT</name></connection>
<intersection>716.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>716.5,2327.5,716.5,2378</points>
<intersection>2327.5 12</intersection>
<intersection>2332.5 13</intersection>
<intersection>2337.5 14</intersection>
<intersection>2342.5 15</intersection>
<intersection>2347.5 16</intersection>
<intersection>2352.5 17</intersection>
<intersection>2357.5 18</intersection>
<intersection>2362.5 19</intersection>
<intersection>2378 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>707.5,2327.5,716.5,2327.5</points>
<connection>
<GID>691</GID>
<name>SEL_0</name></connection>
<intersection>716.5 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>707.5,2332.5,716.5,2332.5</points>
<connection>
<GID>690</GID>
<name>SEL_0</name></connection>
<intersection>716.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>707.5,2337.5,716.5,2337.5</points>
<connection>
<GID>689</GID>
<name>SEL_0</name></connection>
<intersection>716.5 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>707.5,2342.5,716.5,2342.5</points>
<connection>
<GID>692</GID>
<name>SEL_0</name></connection>
<intersection>716.5 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>707.5,2347.5,716.5,2347.5</points>
<connection>
<GID>688</GID>
<name>SEL_0</name></connection>
<intersection>716.5 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>707.5,2352.5,716.5,2352.5</points>
<connection>
<GID>687</GID>
<name>SEL_0</name></connection>
<intersection>716.5 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>707.5,2357.5,716.5,2357.5</points>
<connection>
<GID>686</GID>
<name>SEL_0</name></connection>
<intersection>716.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>707.5,2362.5,716.5,2362.5</points>
<connection>
<GID>675</GID>
<name>SEL_0</name></connection>
<intersection>716.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>891</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>588.5,2355.5,588.5,2359</points>
<connection>
<GID>682</GID>
<name>OUT_1</name></connection>
<intersection>2355.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>588.5,2355.5,590,2355.5</points>
<connection>
<GID>873</GID>
<name>IN_0</name></connection>
<intersection>588.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512,2366.5,512,2370</points>
<connection>
<GID>679</GID>
<name>IN_2</name></connection>
<intersection>2370 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,2370,512,2370</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>512 0</intersection></hsegment></shape></wire>
<wire>
<ID>892</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,2358,589.5,2359</points>
<connection>
<GID>682</GID>
<name>OUT_0</name></connection>
<intersection>2358 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>589.5,2358,590,2358</points>
<connection>
<GID>874</GID>
<name>IN_0</name></connection>
<intersection>589.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,2366.5,511,2367.5</points>
<connection>
<GID>679</GID>
<name>IN_3</name></connection>
<intersection>2367.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>510.5,2367.5,511,2367.5</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>511 0</intersection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>705,2380,705.5,2380</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<connection>
<GID>677</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>524,2363.5,526,2363.5</points>
<connection>
<GID>679</GID>
<name>carry_in</name></connection>
<connection>
<GID>680</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>893</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590,2310.5,590,2311.5</points>
<connection>
<GID>860</GID>
<name>OUT_0</name></connection>
<intersection>2310.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>590,2310.5,590.5,2310.5</points>
<connection>
<GID>887</GID>
<name>IN_0</name></connection>
<intersection>590 0</intersection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>705,2378,705.5,2378</points>
<connection>
<GID>595</GID>
<name>IN_1</name></connection>
<connection>
<GID>678</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>894</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>589,2308,589,2311.5</points>
<connection>
<GID>860</GID>
<name>OUT_1</name></connection>
<intersection>2308 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>589,2308,590.5,2308</points>
<connection>
<GID>886</GID>
<name>IN_0</name></connection>
<intersection>589 2</intersection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>705,2376,705.5,2376</points>
<connection>
<GID>595</GID>
<name>IN_2</name></connection>
<connection>
<GID>683</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578,2364,580,2364</points>
<connection>
<GID>681</GID>
<name>carry_in</name></connection>
<connection>
<GID>682</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>895</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>588,2305.5,588,2311.5</points>
<connection>
<GID>860</GID>
<name>OUT_2</name></connection>
<intersection>2305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>588,2305.5,590.5,2305.5</points>
<connection>
<GID>885</GID>
<name>IN_0</name></connection>
<intersection>588 0</intersection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>565,2367,565,2368</points>
<connection>
<GID>681</GID>
<name>IN_3</name></connection>
<intersection>2368 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>564.5,2368,565,2368</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>565 0</intersection></hsegment></shape></wire>
<wire>
<ID>896</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587,2303,587,2311.5</points>
<connection>
<GID>860</GID>
<name>OUT_3</name></connection>
<intersection>2303 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>587,2303,590.5,2303</points>
<connection>
<GID>880</GID>
<name>IN_0</name></connection>
<intersection>587 0</intersection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>566,2367,566,2370.5</points>
<connection>
<GID>681</GID>
<name>IN_2</name></connection>
<intersection>2370.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>564.5,2370.5,566,2370.5</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>566 0</intersection></hsegment></shape></wire>
<wire>
<ID>897</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>572,2300.5,572,2311.5</points>
<connection>
<GID>859</GID>
<name>OUT_0</name></connection>
<intersection>2300.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>572,2300.5,590.5,2300.5</points>
<connection>
<GID>891</GID>
<name>IN_0</name></connection>
<intersection>572 0</intersection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>532,2366.5,532,2385</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<intersection>2385 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,2385,532,2385</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>532 0</intersection></hsegment></shape></wire>
<wire>
<ID>898</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571,2298,571,2311.5</points>
<connection>
<GID>859</GID>
<name>OUT_1</name></connection>
<intersection>2298 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>571,2298,590.5,2298</points>
<connection>
<GID>890</GID>
<name>IN_0</name></connection>
<intersection>571 0</intersection></hsegment></shape></wire>
<wire>
<ID>899</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>570,2295.5,570,2311.5</points>
<connection>
<GID>859</GID>
<name>OUT_2</name></connection>
<intersection>2295.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>570,2295.5,590.5,2295.5</points>
<connection>
<GID>889</GID>
<name>IN_0</name></connection>
<intersection>570 0</intersection></hsegment></shape></wire>
<wire>
<ID>900</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>569,2293,569,2311.5</points>
<connection>
<GID>859</GID>
<name>OUT_3</name></connection>
<intersection>2293 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>569,2293,590.5,2293</points>
<connection>
<GID>888</GID>
<name>IN_0</name></connection>
<intersection>569 0</intersection></hsegment></shape></wire>
<wire>
<ID>901</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>535.5,2357.5,535.5,2358.5</points>
<connection>
<GID>680</GID>
<name>OUT_0</name></connection>
<intersection>2357.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>535.5,2357.5,536,2357.5</points>
<connection>
<GID>895</GID>
<name>IN_0</name></connection>
<intersection>535.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>902</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>534.5,2355,534.5,2358.5</points>
<connection>
<GID>680</GID>
<name>OUT_1</name></connection>
<intersection>2355 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>534.5,2355,536,2355</points>
<connection>
<GID>894</GID>
<name>IN_0</name></connection>
<intersection>534.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>903</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>533.5,2352.5,533.5,2358.5</points>
<connection>
<GID>680</GID>
<name>OUT_2</name></connection>
<intersection>2352.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>533.5,2352.5,536,2352.5</points>
<connection>
<GID>893</GID>
<name>IN_0</name></connection>
<intersection>533.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>904</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>532.5,2350,532.5,2358.5</points>
<connection>
<GID>680</GID>
<name>OUT_3</name></connection>
<intersection>2350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>532.5,2350,536,2350</points>
<connection>
<GID>892</GID>
<name>IN_0</name></connection>
<intersection>532.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>905</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517.5,2347.5,517.5,2358.5</points>
<connection>
<GID>679</GID>
<name>OUT_0</name></connection>
<intersection>2347.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517.5,2347.5,536,2347.5</points>
<connection>
<GID>899</GID>
<name>IN_0</name></connection>
<intersection>517.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>641.5,2333,641.5,2334</points>
<connection>
<GID>752</GID>
<name>OUT_0</name></connection>
<intersection>2333 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>641.5,2333,642,2333</points>
<connection>
<GID>839</GID>
<name>IN_0</name></connection>
<intersection>641.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>906</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516.5,2345,516.5,2358.5</points>
<connection>
<GID>679</GID>
<name>OUT_1</name></connection>
<intersection>2345 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516.5,2345,536,2345</points>
<connection>
<GID>898</GID>
<name>IN_0</name></connection>
<intersection>516.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640.5,2330.5,640.5,2334</points>
<connection>
<GID>752</GID>
<name>OUT_1</name></connection>
<intersection>2330.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>640.5,2330.5,642,2330.5</points>
<connection>
<GID>840</GID>
<name>IN_0</name></connection>
<intersection>640.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639.5,2328,639.5,2334</points>
<connection>
<GID>752</GID>
<name>OUT_2</name></connection>
<intersection>2328 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639.5,2328,642,2328</points>
<connection>
<GID>842</GID>
<name>IN_0</name></connection>
<intersection>639.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>908</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514.5,2340,514.5,2358.5</points>
<connection>
<GID>679</GID>
<name>OUT_3</name></connection>
<intersection>2340 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514.5,2340,536,2340</points>
<connection>
<GID>896</GID>
<name>IN_0</name></connection>
<intersection>514.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>638.5,2325.5,638.5,2334</points>
<connection>
<GID>752</GID>
<name>OUT_3</name></connection>
<intersection>2325.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>638.5,2325.5,642,2325.5</points>
<connection>
<GID>843</GID>
<name>IN_0</name></connection>
<intersection>638.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>909</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515.5,2342.5,515.5,2358.5</points>
<connection>
<GID>679</GID>
<name>OUT_2</name></connection>
<intersection>2342.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,2342.5,536,2342.5</points>
<connection>
<GID>897</GID>
<name>IN_0</name></connection>
<intersection>515.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>623.5,2323,623.5,2334</points>
<connection>
<GID>751</GID>
<name>OUT_0</name></connection>
<intersection>2323 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>623.5,2323,642,2323</points>
<connection>
<GID>816</GID>
<name>IN_0</name></connection>
<intersection>623.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>910</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>536,2309.5,536,2310.5</points>
<connection>
<GID>903</GID>
<name>IN_0</name></connection>
<connection>
<GID>848</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>622.5,2320.5,622.5,2334</points>
<connection>
<GID>751</GID>
<name>OUT_1</name></connection>
<intersection>2320.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>622.5,2320.5,642,2320.5</points>
<connection>
<GID>818</GID>
<name>IN_0</name></connection>
<intersection>622.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>911</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>535,2307,535,2310.5</points>
<connection>
<GID>848</GID>
<name>OUT_1</name></connection>
<intersection>2307 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>535,2307,536,2307</points>
<connection>
<GID>902</GID>
<name>IN_0</name></connection>
<intersection>535 0</intersection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>621.5,2318,621.5,2334</points>
<connection>
<GID>751</GID>
<name>OUT_2</name></connection>
<intersection>2318 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>621.5,2318,642,2318</points>
<connection>
<GID>820</GID>
<name>IN_0</name></connection>
<intersection>621.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>912</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>534,2304.5,534,2310.5</points>
<connection>
<GID>848</GID>
<name>OUT_2</name></connection>
<intersection>2304.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,2304.5,536,2304.5</points>
<connection>
<GID>901</GID>
<name>IN_0</name></connection>
<intersection>534 0</intersection></hsegment></shape></wire>
<wire>
<ID>913</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>533,2302,533,2310.5</points>
<connection>
<GID>848</GID>
<name>OUT_3</name></connection>
<intersection>2302 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>533,2302,536,2302</points>
<connection>
<GID>900</GID>
<name>IN_0</name></connection>
<intersection>533 0</intersection></hsegment></shape></wire>
<wire>
<ID>914</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>518,2299.5,518,2310.5</points>
<connection>
<GID>847</GID>
<name>OUT_0</name></connection>
<intersection>2299.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>518,2299.5,536,2299.5</points>
<connection>
<GID>907</GID>
<name>IN_0</name></connection>
<intersection>518 0</intersection></hsegment></shape></wire>
<wire>
<ID>915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517,2297,517,2310.5</points>
<connection>
<GID>847</GID>
<name>OUT_1</name></connection>
<intersection>2297 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517,2297,536,2297</points>
<connection>
<GID>906</GID>
<name>IN_0</name></connection>
<intersection>517 0</intersection></hsegment></shape></wire>
<wire>
<ID>916</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516,2294.5,516,2310.5</points>
<connection>
<GID>847</GID>
<name>OUT_2</name></connection>
<intersection>2294.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516,2294.5,536,2294.5</points>
<connection>
<GID>905</GID>
<name>IN_0</name></connection>
<intersection>516 0</intersection></hsegment></shape></wire>
<wire>
<ID>917</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515,2292,515,2310.5</points>
<connection>
<GID>847</GID>
<name>OUT_3</name></connection>
<intersection>2292 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515,2292,536,2292</points>
<connection>
<GID>904</GID>
<name>IN_0</name></connection>
<intersection>515 0</intersection></hsegment></shape></wire>
<wire>
<ID>932</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>649.5,2337.5,649.5,2339</points>
<connection>
<GID>879</GID>
<name>OUT_0</name></connection>
<intersection>2339 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>648,2339,649.5,2339</points>
<connection>
<GID>752</GID>
<name>carry_in</name></connection>
<intersection>649.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>933</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>543,2363.5,543,2365</points>
<connection>
<GID>846</GID>
<name>OUT_0</name></connection>
<intersection>2363.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>542,2363.5,543,2363.5</points>
<connection>
<GID>680</GID>
<name>carry_in</name></connection>
<intersection>543 0</intersection></hsegment></shape></wire>
<wire>
<ID>934</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596.5,2364,596.5,2368</points>
<connection>
<GID>857</GID>
<name>OUT_0</name></connection>
<intersection>2364 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>596,2364,596.5,2364</points>
<connection>
<GID>682</GID>
<name>carry_in</name></connection>
<intersection>596.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>935</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>707.5,2367.5,707.5,2370.5</points>
<connection>
<GID>673</GID>
<name>OUT_0</name></connection>
<intersection>2367.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>706,2367.5,707.5,2367.5</points>
<connection>
<GID>626</GID>
<name>carry_in</name></connection>
<intersection>707.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>937</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>612.5,2332,612.5,2339</points>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>2339 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>612.5,2339,614,2339</points>
<connection>
<GID>751</GID>
<name>carry_out</name></connection>
<intersection>612.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>938</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505,2354,505,2363.5</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>2363.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>505,2363.5,508,2363.5</points>
<connection>
<GID>679</GID>
<name>carry_out</name></connection>
<intersection>505 0</intersection></hsegment></shape></wire>
<wire>
<ID>939</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507,2308,507,2315.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>2315.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>507,2315.5,508.5,2315.5</points>
<connection>
<GID>847</GID>
<name>carry_out</name></connection>
<intersection>507 0</intersection></hsegment></shape></wire>
<wire>
<ID>940</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>559.5,2307.5,559.5,2316.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>2316.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>559.5,2316.5,562.5,2316.5</points>
<connection>
<GID>859</GID>
<name>carry_out</name></connection>
<intersection>559.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>941</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>560,2354.5,560,2364</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>2364 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>560,2364,562,2364</points>
<connection>
<GID>681</GID>
<name>carry_out</name></connection>
<intersection>560 0</intersection></hsegment></shape></wire>
<wire>
<ID>749</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>620.5,2315.5,620.5,2334</points>
<connection>
<GID>751</GID>
<name>OUT_3</name></connection>
<intersection>2315.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>620.5,2315.5,642,2315.5</points>
<connection>
<GID>821</GID>
<name>IN_0</name></connection>
<intersection>620.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>750</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512.5,2318.5,512.5,2322</points>
<connection>
<GID>847</GID>
<name>IN_2</name></connection>
<intersection>2322 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>511,2322,512.5,2322</points>
<connection>
<GID>852</GID>
<name>IN_0</name></connection>
<intersection>512.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>751</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,2318.5,511.5,2319.5</points>
<connection>
<GID>847</GID>
<name>IN_3</name></connection>
<intersection>2319.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>511,2319.5,511.5,2319.5</points>
<connection>
<GID>853</GID>
<name>IN_0</name></connection>
<intersection>511.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>752</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>524.5,2315.5,526.5,2315.5</points>
<connection>
<GID>847</GID>
<name>carry_in</name></connection>
<connection>
<GID>848</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>753</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>532.5,2318.5,532.5,2337</points>
<connection>
<GID>848</GID>
<name>IN_0</name></connection>
<intersection>2337 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,2337,532.5,2337</points>
<connection>
<GID>854</GID>
<name>IN_0</name></connection>
<intersection>532.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>754</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>531.5,2318.5,531.5,2334.5</points>
<connection>
<GID>848</GID>
<name>IN_1</name></connection>
<intersection>2334.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,2334.5,531.5,2334.5</points>
<connection>
<GID>855</GID>
<name>IN_0</name></connection>
<intersection>531.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>755</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530.5,2318.5,530.5,2332</points>
<connection>
<GID>848</GID>
<name>IN_2</name></connection>
<intersection>2332 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,2332,530.5,2332</points>
<connection>
<GID>856</GID>
<name>IN_0</name></connection>
<intersection>530.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>756</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>529.5,2318.5,529.5,2329.5</points>
<connection>
<GID>848</GID>
<name>IN_3</name></connection>
<intersection>2329.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,2329.5,529.5,2329.5</points>
<connection>
<GID>849</GID>
<name>IN_0</name></connection>
<intersection>529.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>757</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514.5,2318.5,514.5,2327</points>
<connection>
<GID>847</GID>
<name>IN_0</name></connection>
<intersection>2327 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>511,2327,514.5,2327</points>
<connection>
<GID>850</GID>
<name>IN_0</name></connection>
<intersection>514.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513.5,2318.5,513.5,2324.5</points>
<connection>
<GID>847</GID>
<name>IN_1</name></connection>
<intersection>2324.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>511,2324.5,513.5,2324.5</points>
<connection>
<GID>851</GID>
<name>IN_0</name></connection>
<intersection>513.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>233.346,6642.04,434.404,6539.25</PageViewport>
<gate>
<ID>1167</ID>
<type>DE_TO</type>
<position>339,6608.5</position>
<input>
<ID>IN_0</ID>1024 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor2</lparam></gate>
<gate>
<ID>1168</ID>
<type>DE_TO</type>
<position>339,6604</position>
<input>
<ID>IN_0</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor3</lparam></gate>
<gate>
<ID>1169</ID>
<type>DE_TO</type>
<position>339,6599.5</position>
<input>
<ID>IN_0</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor4</lparam></gate>
<gate>
<ID>1170</ID>
<type>DE_TO</type>
<position>339,6595</position>
<input>
<ID>IN_0</ID>1025 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor5</lparam></gate>
<gate>
<ID>1171</ID>
<type>DE_TO</type>
<position>339,6590.5</position>
<input>
<ID>IN_0</ID>1022 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor6</lparam></gate>
<gate>
<ID>1172</ID>
<type>DE_TO</type>
<position>339,6586</position>
<input>
<ID>IN_0</ID>1029 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor7</lparam></gate>
<gate>
<ID>1173</ID>
<type>DE_TO</type>
<position>364.5,6615.5</position>
<input>
<ID>IN_0</ID>1031 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor0</lparam></gate>
<gate>
<ID>1174</ID>
<type>DE_TO</type>
<position>364.5,6611</position>
<input>
<ID>IN_0</ID>1032 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor1</lparam></gate>
<gate>
<ID>1175</ID>
<type>DE_TO</type>
<position>364.5,6606.5</position>
<input>
<ID>IN_0</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor2</lparam></gate>
<gate>
<ID>1176</ID>
<type>DE_TO</type>
<position>364.5,6602</position>
<input>
<ID>IN_0</ID>1037 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor3</lparam></gate>
<gate>
<ID>1177</ID>
<type>DE_TO</type>
<position>364.5,6597.5</position>
<input>
<ID>IN_0</ID>1033 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor4</lparam></gate>
<gate>
<ID>1178</ID>
<type>DE_TO</type>
<position>364.5,6593</position>
<input>
<ID>IN_0</ID>1034 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor5</lparam></gate>
<gate>
<ID>1179</ID>
<type>DE_TO</type>
<position>364.5,6588.5</position>
<input>
<ID>IN_0</ID>1030 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor6</lparam></gate>
<gate>
<ID>1180</ID>
<type>DE_TO</type>
<position>364.5,6584</position>
<input>
<ID>IN_0</ID>1035 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor7</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>283.5,6578</position>
<gparam>LABEL_TEXT NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>BA_NAND2</type>
<position>280,6573</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>274.5,6574</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>274.5,6572</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>287,6573</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand0</lparam></gate>
<gate>
<ID>44</ID>
<type>BA_NAND2</type>
<position>280,6568.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>274.5,6569.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>274.5,6567.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>287,6568.5</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand1</lparam></gate>
<gate>
<ID>48</ID>
<type>BA_NAND2</type>
<position>280,6564</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>DA_FROM</type>
<position>274.5,6565</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>274.5,6563</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>287,6564</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand2</lparam></gate>
<gate>
<ID>52</ID>
<type>BA_NAND2</type>
<position>280,6559.5</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>DA_FROM</type>
<position>274.5,6560.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>274.5,6558.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>287,6559.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand3</lparam></gate>
<gate>
<ID>56</ID>
<type>BA_NAND2</type>
<position>280,6555</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>274.5,6556</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>274.5,6554</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>287,6555</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand4</lparam></gate>
<gate>
<ID>60</ID>
<type>BA_NAND2</type>
<position>280,6550.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>91 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>274.5,6551.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>274.5,6549.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>67</ID>
<type>DE_TO</type>
<position>287,6550.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand5</lparam></gate>
<gate>
<ID>71</ID>
<type>BA_NAND2</type>
<position>280,6546</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>274.5,6547</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>274.5,6545</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>75</ID>
<type>DE_TO</type>
<position>287,6546</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand6</lparam></gate>
<gate>
<ID>76</ID>
<type>BA_NAND2</type>
<position>280,6541.5</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>274.5,6542.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>274.5,6540.5</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>80</ID>
<type>DE_TO</type>
<position>287,6541.5</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand7</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>309.5,6578</position>
<gparam>LABEL_TEXT NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>BE_NOR2</type>
<position>308,6573</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>302.5,6574</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>302.5,6572</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>314.5,6573</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor0</lparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>302.5,6567.5</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>87</ID>
<type>DE_TO</type>
<position>314.5,6568.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor1</lparam></gate>
<gate>
<ID>90</ID>
<type>BE_NOR2</type>
<position>308,6568.5</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>DA_FROM</type>
<position>302.5,6569.5</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>302.5,6563</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>98</ID>
<type>DE_TO</type>
<position>314.5,6564</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor2</lparam></gate>
<gate>
<ID>99</ID>
<type>BE_NOR2</type>
<position>308,6564</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>302.5,6565</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>302.5,6558.5</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>314.5,6559.5</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor3</lparam></gate>
<gate>
<ID>103</ID>
<type>BE_NOR2</type>
<position>308,6559.5</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>DA_FROM</type>
<position>302.5,6560.5</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>105</ID>
<type>DA_FROM</type>
<position>302.5,6554</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>314.5,6555</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor4</lparam></gate>
<gate>
<ID>107</ID>
<type>DA_FROM</type>
<position>302.5,6549.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>314.5,6550.5</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor5</lparam></gate>
<gate>
<ID>109</ID>
<type>BE_NOR2</type>
<position>308,6550.5</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>116 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>DA_FROM</type>
<position>302.5,6551.5</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>111</ID>
<type>DA_FROM</type>
<position>302.5,6545</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>112</ID>
<type>DE_TO</type>
<position>314.5,6546</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor6</lparam></gate>
<gate>
<ID>113</ID>
<type>BE_NOR2</type>
<position>308,6546</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>DA_FROM</type>
<position>302.5,6547</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>115</ID>
<type>DA_FROM</type>
<position>302.5,6540.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>116</ID>
<type>DE_TO</type>
<position>314.5,6541.5</position>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor7</lparam></gate>
<gate>
<ID>121</ID>
<type>BE_NOR2</type>
<position>308,6541.5</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>DA_FROM</type>
<position>302.5,6542.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>123</ID>
<type>BE_NOR2</type>
<position>308,6555</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>302.5,6556</position>
<input>
<ID>IN_0</ID>111 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>125</ID>
<type>AE_SMALL_INVERTER</type>
<position>385,6609.5</position>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>380.5,6609.5</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>127</ID>
<type>DE_TO</type>
<position>389.5,6609.5</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx0</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>387,6614</position>
<gparam>LABEL_TEXT NOT</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AE_SMALL_INVERTER</type>
<position>385,6606.5</position>
<input>
<ID>IN_0</ID>128 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>380.5,6606.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>131</ID>
<type>DE_TO</type>
<position>389.5,6606.5</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx1</lparam></gate>
<gate>
<ID>132</ID>
<type>AE_SMALL_INVERTER</type>
<position>385,6603.5</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>380.5,6603.5</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>134</ID>
<type>DE_TO</type>
<position>389.5,6603.5</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx2</lparam></gate>
<gate>
<ID>135</ID>
<type>AE_SMALL_INVERTER</type>
<position>385,6600.5</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>380.5,6600.5</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_TO</type>
<position>389.5,6600.5</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx3</lparam></gate>
<gate>
<ID>139</ID>
<type>AE_SMALL_INVERTER</type>
<position>385,6597.5</position>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>380.5,6597.5</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>141</ID>
<type>DE_TO</type>
<position>389.5,6597.5</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx4</lparam></gate>
<gate>
<ID>142</ID>
<type>AE_SMALL_INVERTER</type>
<position>385,6594.5</position>
<input>
<ID>IN_0</ID>136 </input>
<output>
<ID>OUT_0</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>380.5,6594.5</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_TO</type>
<position>389.5,6594.5</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx5</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_SMALL_INVERTER</type>
<position>385,6591.5</position>
<input>
<ID>IN_0</ID>138 </input>
<output>
<ID>OUT_0</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>146</ID>
<type>DA_FROM</type>
<position>380.5,6591.5</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>147</ID>
<type>DE_TO</type>
<position>389.5,6591.5</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx6</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_SMALL_INVERTER</type>
<position>385,6588.5</position>
<input>
<ID>IN_0</ID>140 </input>
<output>
<ID>OUT_0</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>149</ID>
<type>DA_FROM</type>
<position>380.5,6588.5</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>150</ID>
<type>DE_TO</type>
<position>389.5,6588.5</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx7</lparam></gate>
<gate>
<ID>180</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>340,6556.5</position>
<output>
<ID>A_equal_B</ID>202 </output>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<input>
<ID>IN_2</ID>186 </input>
<input>
<ID>IN_3</ID>185 </input>
<input>
<ID>IN_B_0</ID>189 </input>
<input>
<ID>IN_B_1</ID>190 </input>
<input>
<ID>IN_B_2</ID>191 </input>
<input>
<ID>IN_B_3</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>332.5,6569</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>182</ID>
<type>DA_FROM</type>
<position>332.5,6566.5</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>183</ID>
<type>DA_FROM</type>
<position>332.5,6564</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>332.5,6561.5</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>185</ID>
<type>DA_FROM</type>
<position>377,6569</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>377,6566.5</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>187</ID>
<type>DA_FROM</type>
<position>377,6564</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>188</ID>
<type>DA_FROM</type>
<position>377,6561.5</position>
<input>
<ID>IN_0</ID>193 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>189</ID>
<type>DA_FROM</type>
<position>347.5,6561.5</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>190</ID>
<type>DA_FROM</type>
<position>347.5,6564</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>191</ID>
<type>DA_FROM</type>
<position>347.5,6566.5</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>347.5,6569</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>193</ID>
<type>DA_FROM</type>
<position>392,6569</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>194</ID>
<type>DA_FROM</type>
<position>392,6566.5</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>195</ID>
<type>DA_FROM</type>
<position>392,6564</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>196</ID>
<type>DA_FROM</type>
<position>392,6561.5</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>197</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>384.5,6556.5</position>
<output>
<ID>A_equal_B</ID>203 </output>
<input>
<ID>IN_0</ID>196 </input>
<input>
<ID>IN_1</ID>195 </input>
<input>
<ID>IN_2</ID>194 </input>
<input>
<ID>IN_3</ID>193 </input>
<input>
<ID>IN_B_0</ID>197 </input>
<input>
<ID>IN_B_1</ID>198 </input>
<input>
<ID>IN_B_2</ID>199 </input>
<input>
<ID>IN_B_3</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>198</ID>
<type>DE_TO</type>
<position>364,6565.5</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CMP</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_AND2</type>
<position>361.5,6560</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>361,6574</position>
<gparam>LABEL_TEXT COMPARADOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1029</ID>
<type>AA_LABEL</type>
<position>282,6622</position>
<gparam>LABEL_TEXT AND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1030</ID>
<type>AA_LABEL</type>
<position>309.5,6622.5</position>
<gparam>LABEL_TEXT OR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1031</ID>
<type>AA_LABEL</type>
<position>335,6622.5</position>
<gparam>LABEL_TEXT XOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1032</ID>
<type>AA_LABEL</type>
<position>361,6622.5</position>
<gparam>LABEL_TEXT XNOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1050</ID>
<type>AA_LABEL</type>
<position>325.5,6632</position>
<gparam>LABEL_TEXT Operacoes Portas Logicas</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1052</ID>
<type>AA_LABEL</type>
<position>327,6640.5</position>
<gparam>LABEL_TEXT Unidade logica</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1053</ID>
<type>AA_AND2</type>
<position>281,6617.5</position>
<input>
<ID>IN_0</ID>942 </input>
<input>
<ID>IN_1</ID>943 </input>
<output>
<ID>OUT</ID>1006 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1054</ID>
<type>AA_AND2</type>
<position>281,6613</position>
<input>
<ID>IN_0</ID>944 </input>
<input>
<ID>IN_1</ID>945 </input>
<output>
<ID>OUT</ID>1007 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1055</ID>
<type>AA_AND2</type>
<position>281,6608.5</position>
<input>
<ID>IN_0</ID>957 </input>
<input>
<ID>IN_1</ID>956 </input>
<output>
<ID>OUT</ID>1008 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1056</ID>
<type>AA_AND2</type>
<position>281,6604</position>
<input>
<ID>IN_0</ID>955 </input>
<input>
<ID>IN_1</ID>954 </input>
<output>
<ID>OUT</ID>1009 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1057</ID>
<type>AA_AND2</type>
<position>281,6599.5</position>
<input>
<ID>IN_0</ID>953 </input>
<input>
<ID>IN_1</ID>952 </input>
<output>
<ID>OUT</ID>1010 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1058</ID>
<type>AA_AND2</type>
<position>281,6595</position>
<input>
<ID>IN_0</ID>951 </input>
<input>
<ID>IN_1</ID>950 </input>
<output>
<ID>OUT</ID>1011 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1059</ID>
<type>AA_AND2</type>
<position>281,6590.5</position>
<input>
<ID>IN_0</ID>949 </input>
<input>
<ID>IN_1</ID>948 </input>
<output>
<ID>OUT</ID>1012 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1060</ID>
<type>AA_AND2</type>
<position>281,6586</position>
<input>
<ID>IN_0</ID>947 </input>
<input>
<ID>IN_1</ID>946 </input>
<output>
<ID>OUT</ID>1013 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1061</ID>
<type>AE_OR2</type>
<position>309,6617.5</position>
<input>
<ID>IN_0</ID>960 </input>
<input>
<ID>IN_1</ID>961 </input>
<output>
<ID>OUT</ID>1016 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1062</ID>
<type>AE_OR2</type>
<position>309,6613</position>
<input>
<ID>IN_0</ID>962 </input>
<input>
<ID>IN_1</ID>963 </input>
<output>
<ID>OUT</ID>1015 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1063</ID>
<type>AE_OR2</type>
<position>309,6608.5</position>
<input>
<ID>IN_0</ID>970 </input>
<input>
<ID>IN_1</ID>971 </input>
<output>
<ID>OUT</ID>1014 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1064</ID>
<type>AE_OR2</type>
<position>309,6604</position>
<input>
<ID>IN_0</ID>969 </input>
<input>
<ID>IN_1</ID>968 </input>
<output>
<ID>OUT</ID>1017 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1065</ID>
<type>AE_OR2</type>
<position>309,6599.5</position>
<input>
<ID>IN_0</ID>966 </input>
<input>
<ID>IN_1</ID>967 </input>
<output>
<ID>OUT</ID>1018 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1066</ID>
<type>AE_OR2</type>
<position>309,6595</position>
<input>
<ID>IN_0</ID>964 </input>
<input>
<ID>IN_1</ID>965 </input>
<output>
<ID>OUT</ID>1019 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1067</ID>
<type>AE_OR2</type>
<position>309,6590.5</position>
<input>
<ID>IN_0</ID>972 </input>
<input>
<ID>IN_1</ID>973 </input>
<output>
<ID>OUT</ID>1021 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1068</ID>
<type>AE_OR2</type>
<position>309,6586</position>
<input>
<ID>IN_0</ID>958 </input>
<input>
<ID>IN_1</ID>959 </input>
<output>
<ID>OUT</ID>1020 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1069</ID>
<type>AI_XOR2</type>
<position>333,6617.5</position>
<input>
<ID>IN_0</ID>982 </input>
<input>
<ID>IN_1</ID>983 </input>
<output>
<ID>OUT</ID>1023 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1070</ID>
<type>AI_XOR2</type>
<position>333,6613</position>
<input>
<ID>IN_0</ID>974 </input>
<input>
<ID>IN_1</ID>975 </input>
<output>
<ID>OUT</ID>1026 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1071</ID>
<type>AI_XOR2</type>
<position>333,6608.5</position>
<input>
<ID>IN_0</ID>977 </input>
<input>
<ID>IN_1</ID>976 </input>
<output>
<ID>OUT</ID>1024 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1072</ID>
<type>AI_XOR2</type>
<position>333,6604</position>
<input>
<ID>IN_0</ID>979 </input>
<input>
<ID>IN_1</ID>978 </input>
<output>
<ID>OUT</ID>1027 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1073</ID>
<type>AI_XOR2</type>
<position>333,6599.5</position>
<input>
<ID>IN_0</ID>980 </input>
<input>
<ID>IN_1</ID>981 </input>
<output>
<ID>OUT</ID>1028 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1074</ID>
<type>AI_XOR2</type>
<position>333,6595</position>
<input>
<ID>IN_0</ID>985 </input>
<input>
<ID>IN_1</ID>984 </input>
<output>
<ID>OUT</ID>1025 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1075</ID>
<type>AI_XOR2</type>
<position>333,6590.5</position>
<input>
<ID>IN_0</ID>987 </input>
<input>
<ID>IN_1</ID>986 </input>
<output>
<ID>OUT</ID>1022 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1076</ID>
<type>AI_XOR2</type>
<position>333,6586</position>
<input>
<ID>IN_0</ID>989 </input>
<input>
<ID>IN_1</ID>988 </input>
<output>
<ID>OUT</ID>1029 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1077</ID>
<type>AO_XNOR2</type>
<position>358.5,6615.5</position>
<input>
<ID>IN_0</ID>1002 </input>
<input>
<ID>IN_1</ID>1003 </input>
<output>
<ID>OUT</ID>1031 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1078</ID>
<type>AO_XNOR2</type>
<position>358.5,6611</position>
<input>
<ID>IN_0</ID>1005 </input>
<input>
<ID>IN_1</ID>1004 </input>
<output>
<ID>OUT</ID>1032 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1079</ID>
<type>AO_XNOR2</type>
<position>358.5,6606.5</position>
<input>
<ID>IN_0</ID>990 </input>
<input>
<ID>IN_1</ID>991 </input>
<output>
<ID>OUT</ID>1036 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1080</ID>
<type>AO_XNOR2</type>
<position>358.5,6602</position>
<input>
<ID>IN_0</ID>993 </input>
<input>
<ID>IN_1</ID>992 </input>
<output>
<ID>OUT</ID>1037 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1081</ID>
<type>AO_XNOR2</type>
<position>358.5,6597.5</position>
<input>
<ID>IN_0</ID>996 </input>
<input>
<ID>IN_1</ID>997 </input>
<output>
<ID>OUT</ID>1033 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1082</ID>
<type>AO_XNOR2</type>
<position>358.5,6593</position>
<input>
<ID>IN_0</ID>994 </input>
<input>
<ID>IN_1</ID>995 </input>
<output>
<ID>OUT</ID>1034 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1083</ID>
<type>AO_XNOR2</type>
<position>358.5,6588.5</position>
<input>
<ID>IN_0</ID>998 </input>
<input>
<ID>IN_1</ID>999 </input>
<output>
<ID>OUT</ID>1030 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1084</ID>
<type>AO_XNOR2</type>
<position>358.5,6584</position>
<input>
<ID>IN_0</ID>1001 </input>
<input>
<ID>IN_1</ID>1000 </input>
<output>
<ID>OUT</ID>1035 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1085</ID>
<type>DA_FROM</type>
<position>275,6618.5</position>
<input>
<ID>IN_0</ID>942 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>1086</ID>
<type>DA_FROM</type>
<position>275,6616.5</position>
<input>
<ID>IN_0</ID>943 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>1087</ID>
<type>DA_FROM</type>
<position>275,6614</position>
<input>
<ID>IN_0</ID>944 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>1088</ID>
<type>DA_FROM</type>
<position>275,6612</position>
<input>
<ID>IN_0</ID>945 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>1089</ID>
<type>DA_FROM</type>
<position>275,6609.5</position>
<input>
<ID>IN_0</ID>957 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>1090</ID>
<type>DA_FROM</type>
<position>275,6607.5</position>
<input>
<ID>IN_0</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>1091</ID>
<type>DA_FROM</type>
<position>275,6605</position>
<input>
<ID>IN_0</ID>955 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>1092</ID>
<type>DA_FROM</type>
<position>275,6603</position>
<input>
<ID>IN_0</ID>954 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>1093</ID>
<type>DA_FROM</type>
<position>275,6600.5</position>
<input>
<ID>IN_0</ID>953 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>1094</ID>
<type>DA_FROM</type>
<position>275,6598.5</position>
<input>
<ID>IN_0</ID>952 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>1095</ID>
<type>DA_FROM</type>
<position>275,6596</position>
<input>
<ID>IN_0</ID>951 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>1096</ID>
<type>DA_FROM</type>
<position>275,6594</position>
<input>
<ID>IN_0</ID>950 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>1097</ID>
<type>DA_FROM</type>
<position>275,6591.5</position>
<input>
<ID>IN_0</ID>949 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>1098</ID>
<type>DA_FROM</type>
<position>275,6589.5</position>
<input>
<ID>IN_0</ID>948 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>1099</ID>
<type>DA_FROM</type>
<position>275,6587</position>
<input>
<ID>IN_0</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>1100</ID>
<type>DA_FROM</type>
<position>275,6585</position>
<input>
<ID>IN_0</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>1101</ID>
<type>DA_FROM</type>
<position>303,6618.5</position>
<input>
<ID>IN_0</ID>960 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>1102</ID>
<type>DA_FROM</type>
<position>303,6616.5</position>
<input>
<ID>IN_0</ID>961 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>1103</ID>
<type>DA_FROM</type>
<position>303,6614</position>
<input>
<ID>IN_0</ID>962 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>1104</ID>
<type>DA_FROM</type>
<position>303,6612</position>
<input>
<ID>IN_0</ID>963 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>1105</ID>
<type>DA_FROM</type>
<position>303,6609.5</position>
<input>
<ID>IN_0</ID>970 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>1106</ID>
<type>DA_FROM</type>
<position>303,6607.5</position>
<input>
<ID>IN_0</ID>971 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>1107</ID>
<type>DA_FROM</type>
<position>303,6605</position>
<input>
<ID>IN_0</ID>969 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>1108</ID>
<type>DA_FROM</type>
<position>303,6603</position>
<input>
<ID>IN_0</ID>968 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>1109</ID>
<type>DA_FROM</type>
<position>303,6600.5</position>
<input>
<ID>IN_0</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>1110</ID>
<type>DA_FROM</type>
<position>303,6598.5</position>
<input>
<ID>IN_0</ID>967 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>1111</ID>
<type>DA_FROM</type>
<position>303,6596</position>
<input>
<ID>IN_0</ID>964 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>1112</ID>
<type>DA_FROM</type>
<position>303,6594</position>
<input>
<ID>IN_0</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>1113</ID>
<type>DA_FROM</type>
<position>303,6591.5</position>
<input>
<ID>IN_0</ID>972 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>1114</ID>
<type>DA_FROM</type>
<position>303,6589.5</position>
<input>
<ID>IN_0</ID>973 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>1115</ID>
<type>DA_FROM</type>
<position>303,6587</position>
<input>
<ID>IN_0</ID>958 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>1116</ID>
<type>DA_FROM</type>
<position>303,6585</position>
<input>
<ID>IN_0</ID>959 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>1117</ID>
<type>DA_FROM</type>
<position>327,6618.5</position>
<input>
<ID>IN_0</ID>982 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>1118</ID>
<type>DA_FROM</type>
<position>327,6616.5</position>
<input>
<ID>IN_0</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>1119</ID>
<type>DA_FROM</type>
<position>327,6614</position>
<input>
<ID>IN_0</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>1120</ID>
<type>DA_FROM</type>
<position>327,6612</position>
<input>
<ID>IN_0</ID>975 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>1121</ID>
<type>DA_FROM</type>
<position>327,6609.5</position>
<input>
<ID>IN_0</ID>977 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>1122</ID>
<type>DA_FROM</type>
<position>327,6607.5</position>
<input>
<ID>IN_0</ID>976 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>1123</ID>
<type>DA_FROM</type>
<position>327,6605</position>
<input>
<ID>IN_0</ID>979 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>1124</ID>
<type>DA_FROM</type>
<position>327,6603</position>
<input>
<ID>IN_0</ID>978 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>1125</ID>
<type>DA_FROM</type>
<position>327,6600.5</position>
<input>
<ID>IN_0</ID>980 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>1126</ID>
<type>DA_FROM</type>
<position>327,6598.5</position>
<input>
<ID>IN_0</ID>981 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>1127</ID>
<type>DA_FROM</type>
<position>327,6596</position>
<input>
<ID>IN_0</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>1128</ID>
<type>DA_FROM</type>
<position>327,6594</position>
<input>
<ID>IN_0</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>1129</ID>
<type>DA_FROM</type>
<position>327,6591.5</position>
<input>
<ID>IN_0</ID>987 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>1130</ID>
<type>DA_FROM</type>
<position>327,6589.5</position>
<input>
<ID>IN_0</ID>986 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>1131</ID>
<type>DA_FROM</type>
<position>327,6587</position>
<input>
<ID>IN_0</ID>989 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>1132</ID>
<type>DA_FROM</type>
<position>327,6585</position>
<input>
<ID>IN_0</ID>988 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>1133</ID>
<type>DA_FROM</type>
<position>352.5,6616.5</position>
<input>
<ID>IN_0</ID>1002 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>1134</ID>
<type>DA_FROM</type>
<position>352.5,6614.5</position>
<input>
<ID>IN_0</ID>1003 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>1135</ID>
<type>DA_FROM</type>
<position>352.5,6612</position>
<input>
<ID>IN_0</ID>1005 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>1136</ID>
<type>DA_FROM</type>
<position>352.5,6610</position>
<input>
<ID>IN_0</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>1137</ID>
<type>DA_FROM</type>
<position>352.5,6607.5</position>
<input>
<ID>IN_0</ID>990 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>1138</ID>
<type>DA_FROM</type>
<position>352.5,6605.5</position>
<input>
<ID>IN_0</ID>991 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>1139</ID>
<type>DA_FROM</type>
<position>352.5,6603</position>
<input>
<ID>IN_0</ID>993 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>1140</ID>
<type>DA_FROM</type>
<position>352.5,6601</position>
<input>
<ID>IN_0</ID>992 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>1141</ID>
<type>DA_FROM</type>
<position>352.5,6598.5</position>
<input>
<ID>IN_0</ID>996 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>1142</ID>
<type>DA_FROM</type>
<position>352.5,6596.5</position>
<input>
<ID>IN_0</ID>997 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>1143</ID>
<type>DA_FROM</type>
<position>352.5,6594</position>
<input>
<ID>IN_0</ID>994 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>1144</ID>
<type>DA_FROM</type>
<position>352.5,6592</position>
<input>
<ID>IN_0</ID>995 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>1145</ID>
<type>DA_FROM</type>
<position>352.5,6589.5</position>
<input>
<ID>IN_0</ID>998 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>1146</ID>
<type>DA_FROM</type>
<position>352.5,6587.5</position>
<input>
<ID>IN_0</ID>999 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>1147</ID>
<type>DA_FROM</type>
<position>352.5,6585</position>
<input>
<ID>IN_0</ID>1001 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>1148</ID>
<type>DA_FROM</type>
<position>352.5,6583</position>
<input>
<ID>IN_0</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>1149</ID>
<type>DE_TO</type>
<position>287,6617.5</position>
<input>
<ID>IN_0</ID>1006 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and0</lparam></gate>
<gate>
<ID>1150</ID>
<type>DE_TO</type>
<position>287,6613</position>
<input>
<ID>IN_0</ID>1007 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and1</lparam></gate>
<gate>
<ID>1151</ID>
<type>DE_TO</type>
<position>287,6608.5</position>
<input>
<ID>IN_0</ID>1008 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and2</lparam></gate>
<gate>
<ID>1152</ID>
<type>DE_TO</type>
<position>287,6604</position>
<input>
<ID>IN_0</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and3</lparam></gate>
<gate>
<ID>1153</ID>
<type>DE_TO</type>
<position>287,6599.5</position>
<input>
<ID>IN_0</ID>1010 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and4</lparam></gate>
<gate>
<ID>1154</ID>
<type>DE_TO</type>
<position>287,6595</position>
<input>
<ID>IN_0</ID>1011 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and5</lparam></gate>
<gate>
<ID>1155</ID>
<type>DE_TO</type>
<position>287,6590.5</position>
<input>
<ID>IN_0</ID>1012 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and6</lparam></gate>
<gate>
<ID>1156</ID>
<type>DE_TO</type>
<position>287,6586</position>
<input>
<ID>IN_0</ID>1013 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and7</lparam></gate>
<gate>
<ID>1157</ID>
<type>DE_TO</type>
<position>315,6617.5</position>
<input>
<ID>IN_0</ID>1016 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or0</lparam></gate>
<gate>
<ID>1158</ID>
<type>DE_TO</type>
<position>315,6613</position>
<input>
<ID>IN_0</ID>1015 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or1</lparam></gate>
<gate>
<ID>1159</ID>
<type>DE_TO</type>
<position>315,6608.5</position>
<input>
<ID>IN_0</ID>1014 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or2</lparam></gate>
<gate>
<ID>1160</ID>
<type>DE_TO</type>
<position>315,6604</position>
<input>
<ID>IN_0</ID>1017 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or3</lparam></gate>
<gate>
<ID>1161</ID>
<type>DE_TO</type>
<position>315,6599.5</position>
<input>
<ID>IN_0</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or4</lparam></gate>
<gate>
<ID>1162</ID>
<type>DE_TO</type>
<position>315,6595</position>
<input>
<ID>IN_0</ID>1019 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or5</lparam></gate>
<gate>
<ID>1163</ID>
<type>DE_TO</type>
<position>315,6590.5</position>
<input>
<ID>IN_0</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or6</lparam></gate>
<gate>
<ID>1164</ID>
<type>DE_TO</type>
<position>315,6586</position>
<input>
<ID>IN_0</ID>1020 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or7</lparam></gate>
<gate>
<ID>1165</ID>
<type>DE_TO</type>
<position>339,6617.5</position>
<input>
<ID>IN_0</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor0</lparam></gate>
<gate>
<ID>1166</ID>
<type>DE_TO</type>
<position>339,6613</position>
<input>
<ID>IN_0</ID>1026 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor1</lparam></gate>
<wire>
<ID>965</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6594,306,6594</points>
<connection>
<GID>1112</GID>
<name>IN_0</name></connection>
<connection>
<GID>1066</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379.5,6560.5,379.5,6561.5</points>
<connection>
<GID>197</GID>
<name>IN_3</name></connection>
<intersection>6561.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,6561.5,379.5,6561.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>379.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>966</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6600.5,306,6600.5</points>
<connection>
<GID>1109</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380.5,6560.5,380.5,6564</points>
<connection>
<GID>197</GID>
<name>IN_2</name></connection>
<intersection>6564 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,6564,380.5,6564</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>380.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>967</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6598.5,306,6598.5</points>
<connection>
<GID>1110</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381.5,6560.5,381.5,6566.5</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>6566.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,6566.5,381.5,6566.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>381.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>968</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6603,306,6603</points>
<connection>
<GID>1108</GID>
<name>IN_0</name></connection>
<connection>
<GID>1064</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382.5,6560.5,382.5,6569</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>6569 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,6569,382.5,6569</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>382.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>969</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6605,306,6605</points>
<connection>
<GID>1107</GID>
<name>IN_0</name></connection>
<connection>
<GID>1064</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389.5,6560.5,389.5,6561.5</points>
<connection>
<GID>197</GID>
<name>IN_B_0</name></connection>
<intersection>6561.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>389.5,6561.5,390,6561.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>389.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>970</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6609.5,306,6609.5</points>
<connection>
<GID>1105</GID>
<name>IN_0</name></connection>
<connection>
<GID>1063</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388.5,6560.5,388.5,6564</points>
<connection>
<GID>197</GID>
<name>IN_B_1</name></connection>
<intersection>6564 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>388.5,6564,390,6564</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>388.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>971</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6607.5,306,6607.5</points>
<connection>
<GID>1106</GID>
<name>IN_0</name></connection>
<connection>
<GID>1063</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>387.5,6560.5,387.5,6566.5</points>
<connection>
<GID>197</GID>
<name>IN_B_2</name></connection>
<intersection>6566.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>387.5,6566.5,390,6566.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>387.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>972</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6591.5,306,6591.5</points>
<connection>
<GID>1113</GID>
<name>IN_0</name></connection>
<connection>
<GID>1067</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>386.5,6560.5,386.5,6569</points>
<connection>
<GID>197</GID>
<name>IN_B_3</name></connection>
<intersection>6569 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>386.5,6569,390,6569</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>386.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>973</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6589.5,306,6589.5</points>
<connection>
<GID>1114</GID>
<name>IN_0</name></connection>
<connection>
<GID>1067</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,6563,361.5,6565.5</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<intersection>6565.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361.5,6565.5,362,6565.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>361.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>974</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329,6614,330,6614</points>
<connection>
<GID>1119</GID>
<name>IN_0</name></connection>
<connection>
<GID>1070</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>360.5,6552.5,360.5,6557</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>6552.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>331,6552.5,360.5,6552.5</points>
<intersection>331 2</intersection>
<intersection>360.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>331,6552.5,331,6556.5</points>
<intersection>6552.5 1</intersection>
<intersection>6556.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>331,6556.5,332,6556.5</points>
<connection>
<GID>180</GID>
<name>A_equal_B</name></connection>
<intersection>331 2</intersection></hsegment></shape></wire>
<wire>
<ID>975</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329,6612,330,6612</points>
<connection>
<GID>1120</GID>
<name>IN_0</name></connection>
<connection>
<GID>1070</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362.5,6556.5,362.5,6557</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>6556.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362.5,6556.5,376.5,6556.5</points>
<connection>
<GID>197</GID>
<name>A_equal_B</name></connection>
<intersection>362.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>976</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6607.5,330,6607.5</points>
<connection>
<GID>1122</GID>
<name>IN_0</name></connection>
<connection>
<GID>1071</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>977</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329,6609.5,330,6609.5</points>
<connection>
<GID>1121</GID>
<name>IN_0</name></connection>
<connection>
<GID>1071</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>978</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6603,330,6603</points>
<connection>
<GID>1124</GID>
<name>IN_0</name></connection>
<connection>
<GID>1072</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>979</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6605,330,6605</points>
<connection>
<GID>1123</GID>
<name>IN_0</name></connection>
<connection>
<GID>1072</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>980</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6600.5,330,6600.5</points>
<connection>
<GID>1125</GID>
<name>IN_0</name></connection>
<connection>
<GID>1073</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>981</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6598.5,330,6598.5</points>
<connection>
<GID>1126</GID>
<name>IN_0</name></connection>
<connection>
<GID>1073</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>982</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329,6618.5,330,6618.5</points>
<connection>
<GID>1117</GID>
<name>IN_0</name></connection>
<connection>
<GID>1069</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>983</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329,6616.5,330,6616.5</points>
<connection>
<GID>1118</GID>
<name>IN_0</name></connection>
<connection>
<GID>1069</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>984</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6594,330,6594</points>
<connection>
<GID>1128</GID>
<name>IN_0</name></connection>
<connection>
<GID>1074</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>985</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6596,330,6596</points>
<connection>
<GID>1127</GID>
<name>IN_0</name></connection>
<connection>
<GID>1074</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>986</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6589.5,330,6589.5</points>
<connection>
<GID>1130</GID>
<name>IN_0</name></connection>
<connection>
<GID>1075</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>987</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6591.5,330,6591.5</points>
<connection>
<GID>1129</GID>
<name>IN_0</name></connection>
<connection>
<GID>1075</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>988</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6585,330,6585</points>
<connection>
<GID>1132</GID>
<name>IN_0</name></connection>
<connection>
<GID>1076</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>989</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>329,6587,330,6587</points>
<connection>
<GID>1131</GID>
<name>IN_0</name></connection>
<connection>
<GID>1076</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>990</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6607.5,355.5,6607.5</points>
<connection>
<GID>1079</GID>
<name>IN_0</name></connection>
<connection>
<GID>1137</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>991</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6605.5,355.5,6605.5</points>
<connection>
<GID>1079</GID>
<name>IN_1</name></connection>
<connection>
<GID>1138</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>992</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6601,355.5,6601</points>
<connection>
<GID>1080</GID>
<name>IN_1</name></connection>
<connection>
<GID>1140</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>993</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6603,355.5,6603</points>
<connection>
<GID>1080</GID>
<name>IN_0</name></connection>
<connection>
<GID>1139</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>994</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6594,355.5,6594</points>
<connection>
<GID>1082</GID>
<name>IN_0</name></connection>
<connection>
<GID>1143</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>995</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6592,355.5,6592</points>
<connection>
<GID>1082</GID>
<name>IN_1</name></connection>
<connection>
<GID>1144</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>996</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6598.5,355.5,6598.5</points>
<connection>
<GID>1081</GID>
<name>IN_0</name></connection>
<connection>
<GID>1141</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>997</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6596.5,355.5,6596.5</points>
<connection>
<GID>1081</GID>
<name>IN_1</name></connection>
<connection>
<GID>1142</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>998</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6589.5,355.5,6589.5</points>
<connection>
<GID>1083</GID>
<name>IN_0</name></connection>
<connection>
<GID>1145</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>999</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6587.5,355.5,6587.5</points>
<connection>
<GID>1083</GID>
<name>IN_1</name></connection>
<connection>
<GID>1146</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1000</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6583,355.5,6583</points>
<connection>
<GID>1084</GID>
<name>IN_1</name></connection>
<connection>
<GID>1148</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1001</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6585,355.5,6585</points>
<connection>
<GID>1084</GID>
<name>IN_0</name></connection>
<connection>
<GID>1147</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1002</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6616.5,355.5,6616.5</points>
<connection>
<GID>1077</GID>
<name>IN_0</name></connection>
<connection>
<GID>1133</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1003</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6614.5,355.5,6614.5</points>
<connection>
<GID>1077</GID>
<name>IN_1</name></connection>
<connection>
<GID>1134</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1004</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6610,355.5,6610</points>
<connection>
<GID>1078</GID>
<name>IN_1</name></connection>
<connection>
<GID>1136</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1005</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>354.5,6612,355.5,6612</points>
<connection>
<GID>1078</GID>
<name>IN_0</name></connection>
<connection>
<GID>1135</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1006</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>284,6617.5,285,6617.5</points>
<connection>
<GID>1149</GID>
<name>IN_0</name></connection>
<connection>
<GID>1053</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1007</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>284,6613,285,6613</points>
<connection>
<GID>1150</GID>
<name>IN_0</name></connection>
<connection>
<GID>1054</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1008</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>284,6608.5,285,6608.5</points>
<connection>
<GID>1151</GID>
<name>IN_0</name></connection>
<connection>
<GID>1055</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1009</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>284,6604,285,6604</points>
<connection>
<GID>1152</GID>
<name>IN_0</name></connection>
<connection>
<GID>1056</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1010</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>284,6599.5,285,6599.5</points>
<connection>
<GID>1153</GID>
<name>IN_0</name></connection>
<connection>
<GID>1057</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1011</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>284,6595,285,6595</points>
<connection>
<GID>1154</GID>
<name>IN_0</name></connection>
<connection>
<GID>1058</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1012</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>284,6590.5,285,6590.5</points>
<connection>
<GID>1155</GID>
<name>IN_0</name></connection>
<connection>
<GID>1059</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1013</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>284,6586,285,6586</points>
<connection>
<GID>1156</GID>
<name>IN_0</name></connection>
<connection>
<GID>1060</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1014</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>312,6608.5,313,6608.5</points>
<connection>
<GID>1159</GID>
<name>IN_0</name></connection>
<connection>
<GID>1063</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1015</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>312,6613,313,6613</points>
<connection>
<GID>1158</GID>
<name>IN_0</name></connection>
<connection>
<GID>1062</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1016</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>312,6617.5,313,6617.5</points>
<connection>
<GID>1157</GID>
<name>IN_0</name></connection>
<connection>
<GID>1061</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1017</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>312,6604,313,6604</points>
<connection>
<GID>1160</GID>
<name>IN_0</name></connection>
<connection>
<GID>1064</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1018</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>312,6599.5,313,6599.5</points>
<connection>
<GID>1161</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1019</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>312,6595,313,6595</points>
<connection>
<GID>1162</GID>
<name>IN_0</name></connection>
<connection>
<GID>1066</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1020</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>312,6586,313,6586</points>
<connection>
<GID>1164</GID>
<name>IN_0</name></connection>
<connection>
<GID>1068</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1021</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>312,6590.5,313,6590.5</points>
<connection>
<GID>1163</GID>
<name>IN_0</name></connection>
<connection>
<GID>1067</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1022</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>336,6590.5,337,6590.5</points>
<connection>
<GID>1171</GID>
<name>IN_0</name></connection>
<connection>
<GID>1075</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1023</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>336,6617.5,337,6617.5</points>
<connection>
<GID>1165</GID>
<name>IN_0</name></connection>
<connection>
<GID>1069</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1024</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>336,6608.5,337,6608.5</points>
<connection>
<GID>1167</GID>
<name>IN_0</name></connection>
<connection>
<GID>1071</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1025</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>336,6595,337,6595</points>
<connection>
<GID>1170</GID>
<name>IN_0</name></connection>
<connection>
<GID>1074</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1026</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>336,6613,337,6613</points>
<connection>
<GID>1166</GID>
<name>IN_0</name></connection>
<connection>
<GID>1070</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1027</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>336,6604,337,6604</points>
<connection>
<GID>1168</GID>
<name>IN_0</name></connection>
<connection>
<GID>1072</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1028</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>336,6599.5,337,6599.5</points>
<connection>
<GID>1169</GID>
<name>IN_0</name></connection>
<connection>
<GID>1073</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1029</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>336,6586,337,6586</points>
<connection>
<GID>1172</GID>
<name>IN_0</name></connection>
<connection>
<GID>1076</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1030</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>361.5,6588.5,362.5,6588.5</points>
<connection>
<GID>1083</GID>
<name>OUT</name></connection>
<connection>
<GID>1179</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>361.5,6615.5,362.5,6615.5</points>
<connection>
<GID>1077</GID>
<name>OUT</name></connection>
<connection>
<GID>1173</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1032</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>361.5,6611,362.5,6611</points>
<connection>
<GID>1078</GID>
<name>OUT</name></connection>
<connection>
<GID>1174</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1033</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>361.5,6597.5,362.5,6597.5</points>
<connection>
<GID>1081</GID>
<name>OUT</name></connection>
<connection>
<GID>1177</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>361.5,6593,362.5,6593</points>
<connection>
<GID>1082</GID>
<name>OUT</name></connection>
<connection>
<GID>1178</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>361.5,6584,362.5,6584</points>
<connection>
<GID>1084</GID>
<name>OUT</name></connection>
<connection>
<GID>1180</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>361.5,6606.5,362.5,6606.5</points>
<connection>
<GID>1079</GID>
<name>OUT</name></connection>
<connection>
<GID>1175</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>361.5,6602,362.5,6602</points>
<connection>
<GID>1080</GID>
<name>OUT</name></connection>
<connection>
<GID>1176</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6574,277,6574</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6572,277,6572</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283,6573,285,6573</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6569.5,277,6569.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6567.5,277,6567.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>283,6568.5,285,6568.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6565,277,6565</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6563,277,6563</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283,6564,285,6564</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<connection>
<GID>51</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6560.5,277,6560.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6558.5,277,6558.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<connection>
<GID>54</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283,6559.5,285,6559.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6556,277,6556</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6554,277,6554</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283,6555,285,6555</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6551.5,277,6551.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6549.5,277,6549.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>283,6550.5,285,6550.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6547,277,6547</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6545,277,6545</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283,6546,285,6546</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<connection>
<GID>75</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6542.5,277,6542.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,6540.5,277,6540.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283,6541.5,285,6541.5</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>80</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304.5,6574,305,6574</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<connection>
<GID>83</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304.5,6572,305,6572</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<connection>
<GID>84</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>311,6573,312.5,6573</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<connection>
<GID>85</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304.5,6569.5,305,6569.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>304.5,6567.5,305,6567.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<connection>
<GID>90</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,6568.5,312.5,6568.5</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304.5,6565,305,6565</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>25</ID>
<points>304.5,6563,305,6563</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,6564,312.5,6564</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304.5,6560.5,305,6560.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>104</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>304.5,6558.5,305,6558.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<connection>
<GID>103</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,6559.5,312.5,6559.5</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304.5,6556,305,6556</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<connection>
<GID>124</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>304.5,6554,305,6554</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<connection>
<GID>123</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,6555,312.5,6555</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304.5,6551.5,305,6551.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>304.5,6549.5,305,6549.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<connection>
<GID>109</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,6550.5,312.5,6550.5</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304.5,6547,305,6547</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<connection>
<GID>114</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>25</ID>
<points>304.5,6545,305,6545</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<connection>
<GID>113</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,6546,312.5,6546</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304.5,6542.5,305,6542.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>304.5,6540.5,305,6540.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,6541.5,312.5,6541.5</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<connection>
<GID>116</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,6609.5,383,6609.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>10</ID>
<points>387,6609.5,387.5,6609.5</points>
<connection>
<GID>125</GID>
<name>OUT_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,6606.5,383,6606.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>10</ID>
<points>387,6606.5,387.5,6606.5</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,6603.5,383,6603.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>10</ID>
<points>387,6603.5,387.5,6603.5</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,6600.5,383,6600.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>10</ID>
<points>387,6600.5,387.5,6600.5</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,6597.5,383,6597.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>387,6597.5,387.5,6597.5</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,6594.5,383,6594.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>387,6594.5,387.5,6594.5</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<connection>
<GID>144</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,6591.5,383,6591.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>387,6591.5,387.5,6591.5</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<connection>
<GID>147</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,6588.5,383,6588.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>387,6588.5,387.5,6588.5</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<connection>
<GID>150</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>942</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6618.5,278,6618.5</points>
<connection>
<GID>1085</GID>
<name>IN_0</name></connection>
<connection>
<GID>1053</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>943</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6616.5,278,6616.5</points>
<connection>
<GID>1086</GID>
<name>IN_0</name></connection>
<connection>
<GID>1053</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>944</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6614,278,6614</points>
<connection>
<GID>1087</GID>
<name>IN_0</name></connection>
<connection>
<GID>1054</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>945</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6612,278,6612</points>
<connection>
<GID>1088</GID>
<name>IN_0</name></connection>
<connection>
<GID>1054</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>946</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6585,278,6585</points>
<connection>
<GID>1100</GID>
<name>IN_0</name></connection>
<connection>
<GID>1060</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>947</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6587,278,6587</points>
<connection>
<GID>1099</GID>
<name>IN_0</name></connection>
<connection>
<GID>1060</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>948</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6589.5,278,6589.5</points>
<connection>
<GID>1098</GID>
<name>IN_0</name></connection>
<connection>
<GID>1059</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>949</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6591.5,278,6591.5</points>
<connection>
<GID>1097</GID>
<name>IN_0</name></connection>
<connection>
<GID>1059</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>950</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6594,278,6594</points>
<connection>
<GID>1096</GID>
<name>IN_0</name></connection>
<connection>
<GID>1058</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>951</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6596,278,6596</points>
<connection>
<GID>1095</GID>
<name>IN_0</name></connection>
<connection>
<GID>1058</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>952</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6598.5,278,6598.5</points>
<connection>
<GID>1094</GID>
<name>IN_0</name></connection>
<connection>
<GID>1057</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>953</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6600.5,278,6600.5</points>
<connection>
<GID>1093</GID>
<name>IN_0</name></connection>
<connection>
<GID>1057</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>954</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6603,278,6603</points>
<connection>
<GID>1092</GID>
<name>IN_0</name></connection>
<connection>
<GID>1056</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>955</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6605,278,6605</points>
<connection>
<GID>1091</GID>
<name>IN_0</name></connection>
<connection>
<GID>1056</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>956</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6607.5,278,6607.5</points>
<connection>
<GID>1090</GID>
<name>IN_0</name></connection>
<connection>
<GID>1055</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>957</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,6609.5,278,6609.5</points>
<connection>
<GID>1089</GID>
<name>IN_0</name></connection>
<connection>
<GID>1055</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335,6560.5,335,6561.5</points>
<connection>
<GID>180</GID>
<name>IN_3</name></connection>
<intersection>6561.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>334.5,6561.5,335,6561.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>335 0</intersection></hsegment></shape></wire>
<wire>
<ID>958</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6587,306,6587</points>
<connection>
<GID>1115</GID>
<name>IN_0</name></connection>
<connection>
<GID>1068</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336,6560.5,336,6564</points>
<connection>
<GID>180</GID>
<name>IN_2</name></connection>
<intersection>6564 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334.5,6564,336,6564</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>336 0</intersection></hsegment></shape></wire>
<wire>
<ID>959</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6585,306,6585</points>
<connection>
<GID>1116</GID>
<name>IN_0</name></connection>
<connection>
<GID>1068</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,6560.5,337,6566.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>6566.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334.5,6566.5,337,6566.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>337 0</intersection></hsegment></shape></wire>
<wire>
<ID>960</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6618.5,306,6618.5</points>
<connection>
<GID>1101</GID>
<name>IN_0</name></connection>
<connection>
<GID>1061</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338,6560.5,338,6569</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>6569 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334.5,6569,338,6569</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>338 0</intersection></hsegment></shape></wire>
<wire>
<ID>961</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6616.5,306,6616.5</points>
<connection>
<GID>1102</GID>
<name>IN_0</name></connection>
<connection>
<GID>1061</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345,6560.5,345,6561.5</points>
<connection>
<GID>180</GID>
<name>IN_B_0</name></connection>
<intersection>6561.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345,6561.5,345.5,6561.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>345 0</intersection></hsegment></shape></wire>
<wire>
<ID>962</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6614,306,6614</points>
<connection>
<GID>1103</GID>
<name>IN_0</name></connection>
<connection>
<GID>1062</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344,6560.5,344,6564</points>
<connection>
<GID>180</GID>
<name>IN_B_1</name></connection>
<intersection>6564 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344,6564,345.5,6564</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>344 0</intersection></hsegment></shape></wire>
<wire>
<ID>963</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6612,306,6612</points>
<connection>
<GID>1104</GID>
<name>IN_0</name></connection>
<connection>
<GID>1062</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>343,6560.5,343,6566.5</points>
<connection>
<GID>180</GID>
<name>IN_B_2</name></connection>
<intersection>6566.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>343,6566.5,345.5,6566.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>343 0</intersection></hsegment></shape></wire>
<wire>
<ID>964</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,6596,306,6596</points>
<connection>
<GID>1111</GID>
<name>IN_0</name></connection>
<connection>
<GID>1066</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342,6560.5,342,6569</points>
<connection>
<GID>180</GID>
<name>IN_B_3</name></connection>
<intersection>6569 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,6569,345.5,6569</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>342 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>212.625,6614.02,471.275,6481.79</PageViewport>
<gate>
<ID>1556</ID>
<type>AA_MUX_2x1</type>
<position>393.5,6574.5</position>
<input>
<ID>IN_0</ID>1288 </input>
<input>
<ID>IN_1</ID>1296 </input>
<output>
<ID>OUT</ID>1299 </output>
<input>
<ID>SEL_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1557</ID>
<type>AA_MUX_2x1</type>
<position>393.5,6569.5</position>
<input>
<ID>IN_0</ID>1287 </input>
<input>
<ID>IN_1</ID>1295 </input>
<output>
<ID>OUT</ID>1300 </output>
<input>
<ID>SEL_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1558</ID>
<type>AA_MUX_2x1</type>
<position>393.5,6564.5</position>
<input>
<ID>IN_0</ID>1286 </input>
<input>
<ID>IN_1</ID>1294 </input>
<output>
<ID>OUT</ID>1301 </output>
<input>
<ID>SEL_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1559</ID>
<type>AA_MUX_2x1</type>
<position>393.5,6554.5</position>
<input>
<ID>IN_0</ID>1284 </input>
<input>
<ID>IN_1</ID>1292 </input>
<output>
<ID>OUT</ID>1303 </output>
<input>
<ID>SEL_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1560</ID>
<type>AA_MUX_2x1</type>
<position>393.5,6549.5</position>
<input>
<ID>IN_0</ID>1283 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1304 </output>
<input>
<ID>SEL_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1561</ID>
<type>AA_MUX_2x1</type>
<position>393.5,6544.5</position>
<input>
<ID>IN_0</ID>1282 </input>
<input>
<ID>IN_1</ID>1290 </input>
<output>
<ID>OUT</ID>1305 </output>
<input>
<ID>SEL_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1562</ID>
<type>AA_MUX_2x1</type>
<position>393.5,6559.5</position>
<input>
<ID>IN_0</ID>1285 </input>
<input>
<ID>IN_1</ID>1293 </input>
<output>
<ID>OUT</ID>1302 </output>
<input>
<ID>SEL_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1563</ID>
<type>DA_FROM</type>
<position>389,6563.5</position>
<input>
<ID>IN_0</ID>1286 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa4</lparam></gate>
<gate>
<ID>1564</ID>
<type>DA_FROM</type>
<position>389,6558.5</position>
<input>
<ID>IN_0</ID>1285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa3</lparam></gate>
<gate>
<ID>1565</ID>
<type>DA_FROM</type>
<position>389,6553.5</position>
<input>
<ID>IN_0</ID>1284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa2</lparam></gate>
<gate>
<ID>1566</ID>
<type>DA_FROM</type>
<position>389,6548.5</position>
<input>
<ID>IN_0</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa1</lparam></gate>
<gate>
<ID>1567</ID>
<type>DA_FROM</type>
<position>389,6543.5</position>
<input>
<ID>IN_0</ID>1282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa0</lparam></gate>
<gate>
<ID>1568</ID>
<type>DA_FROM</type>
<position>389,6578.5</position>
<input>
<ID>IN_0</ID>1281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa7</lparam></gate>
<gate>
<ID>1569</ID>
<type>DA_FROM</type>
<position>389,6573.5</position>
<input>
<ID>IN_0</ID>1288 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa6</lparam></gate>
<gate>
<ID>1570</ID>
<type>DA_FROM</type>
<position>389,6568.5</position>
<input>
<ID>IN_0</ID>1287 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa5</lparam></gate>
<gate>
<ID>1571</ID>
<type>DA_FROM</type>
<position>391.5,6584.5</position>
<input>
<ID>IN_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s3</lparam></gate>
<gate>
<ID>1572</ID>
<type>AA_LABEL</type>
<position>424,6596.5</position>
<gparam>LABEL_TEXT Mux 2-1 (*faz a juncao do Mux Aritmetico</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1573</ID>
<type>DA_FROM</type>
<position>389,6545.5</position>
<input>
<ID>IN_0</ID>1290 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol0</lparam></gate>
<gate>
<ID>1574</ID>
<type>DA_FROM</type>
<position>389,6550.5</position>
<input>
<ID>IN_0</ID>1291 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol1</lparam></gate>
<gate>
<ID>1575</ID>
<type>DA_FROM</type>
<position>389,6555.5</position>
<input>
<ID>IN_0</ID>1292 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol2</lparam></gate>
<gate>
<ID>1576</ID>
<type>DA_FROM</type>
<position>389,6560.5</position>
<input>
<ID>IN_0</ID>1293 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol3</lparam></gate>
<gate>
<ID>1577</ID>
<type>DA_FROM</type>
<position>389,6565.5</position>
<input>
<ID>IN_0</ID>1294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol4</lparam></gate>
<gate>
<ID>1578</ID>
<type>DA_FROM</type>
<position>389,6570.5</position>
<input>
<ID>IN_0</ID>1295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol5</lparam></gate>
<gate>
<ID>1579</ID>
<type>DA_FROM</type>
<position>389,6575.5</position>
<input>
<ID>IN_0</ID>1296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol6</lparam></gate>
<gate>
<ID>1580</ID>
<type>DA_FROM</type>
<position>389,6580.5</position>
<input>
<ID>IN_0</ID>1297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol7</lparam></gate>
<gate>
<ID>1582</ID>
<type>AA_LABEL</type>
<position>434,6590.5</position>
<gparam>LABEL_TEXT e</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1584</ID>
<type>AA_LABEL</type>
<position>433,6584</position>
<gparam>LABEL_TEXT  Mux Logico)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1215</ID>
<type>DM_NOR8</type>
<position>423.5,6513.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1122 </input>
<input>
<ID>IN_2</ID>1123 </input>
<input>
<ID>IN_3</ID>1124 </input>
<input>
<ID>IN_4</ID>1101 </input>
<input>
<ID>IN_5</ID>1120 </input>
<input>
<ID>IN_6</ID>1121 </input>
<input>
<ID>IN_7</ID>1125 </input>
<output>
<ID>OUT</ID>1100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1216</ID>
<type>DA_FROM</type>
<position>411,6520.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g0</lparam></gate>
<gate>
<ID>1217</ID>
<type>DA_FROM</type>
<position>411,6518.5</position>
<input>
<ID>IN_0</ID>1122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g1</lparam></gate>
<gate>
<ID>1218</ID>
<type>DA_FROM</type>
<position>411,6514.5</position>
<input>
<ID>IN_0</ID>1124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g3</lparam></gate>
<gate>
<ID>1219</ID>
<type>DA_FROM</type>
<position>411,6510.5</position>
<input>
<ID>IN_0</ID>1121 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g5</lparam></gate>
<gate>
<ID>1220</ID>
<type>DA_FROM</type>
<position>411,6512.5</position>
<input>
<ID>IN_0</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g4</lparam></gate>
<gate>
<ID>1221</ID>
<type>DA_FROM</type>
<position>411,6516.5</position>
<input>
<ID>IN_0</ID>1123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g2</lparam></gate>
<gate>
<ID>1222</ID>
<type>DA_FROM</type>
<position>411,6508.5</position>
<input>
<ID>IN_0</ID>1120 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g6</lparam></gate>
<gate>
<ID>1223</ID>
<type>DA_FROM</type>
<position>411,6506.5</position>
<input>
<ID>IN_0</ID>1101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g7</lparam></gate>
<gate>
<ID>1225</ID>
<type>AI_MUX_8x1</type>
<position>397,6509</position>
<input>
<ID>IN_0</ID>1111 </input>
<input>
<ID>IN_1</ID>1102 </input>
<input>
<ID>IN_2</ID>1103 </input>
<input>
<ID>IN_3</ID>1104 </input>
<input>
<ID>IN_4</ID>1111 </input>
<input>
<ID>IN_5</ID>1105 </input>
<input>
<ID>IN_6</ID>1106 </input>
<input>
<ID>IN_7</ID>1107 </input>
<output>
<ID>OUT</ID>1099 </output>
<input>
<ID>SEL_0</ID>1110 </input>
<input>
<ID>SEL_1</ID>1109 </input>
<input>
<ID>SEL_2</ID>1108 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1226</ID>
<type>AA_LABEL</type>
<position>406,6529.5</position>
<gparam>LABEL_TEXT Unidade de Flags</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>1227</ID>
<type>DE_TO</type>
<position>403.5,6509</position>
<input>
<ID>IN_0</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c</lparam></gate>
<gate>
<ID>1228</ID>
<type>DE_TO</type>
<position>430.5,6513.5</position>
<input>
<ID>IN_0</ID>1100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID z</lparam></gate>
<gate>
<ID>1229</ID>
<type>DA_FROM</type>
<position>386.5,6508.5</position>
<input>
<ID>IN_0</ID>1104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cs</lparam></gate>
<gate>
<ID>1230</ID>
<type>DA_FROM</type>
<position>386.5,6504.5</position>
<input>
<ID>IN_0</ID>1102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cix</lparam></gate>
<gate>
<ID>1231</ID>
<type>DA_FROM</type>
<position>386.5,6506.5</position>
<input>
<ID>IN_0</ID>1103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cdx</lparam></gate>
<gate>
<ID>1232</ID>
<type>DA_FROM</type>
<position>386.5,6512.5</position>
<input>
<ID>IN_0</ID>1106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cdy</lparam></gate>
<gate>
<ID>1233</ID>
<type>DA_FROM</type>
<position>386.5,6510.5</position>
<input>
<ID>IN_0</ID>1105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ciy</lparam></gate>
<gate>
<ID>1234</ID>
<type>DA_FROM</type>
<position>386.5,6514.5</position>
<input>
<ID>IN_0</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cs</lparam></gate>
<gate>
<ID>1235</ID>
<type>DA_FROM</type>
<position>393,6521</position>
<input>
<ID>IN_0</ID>1110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1236</ID>
<type>DA_FROM</type>
<position>393,6517</position>
<input>
<ID>IN_0</ID>1108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1237</ID>
<type>DA_FROM</type>
<position>393,6519</position>
<input>
<ID>IN_0</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1238</ID>
<type>FF_GND</type>
<position>390,6502</position>
<output>
<ID>OUT_0</ID>1111 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1239</ID>
<type>AA_AND2</type>
<position>424,6493</position>
<input>
<ID>IN_0</ID>1114 </input>
<input>
<ID>IN_1</ID>1112 </input>
<output>
<ID>OUT</ID>1118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1240</ID>
<type>DE_TO</type>
<position>394.5,6493</position>
<input>
<ID>IN_0</ID>1097 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID n</lparam></gate>
<gate>
<ID>1241</ID>
<type>AI_XOR2</type>
<position>415.5,6489.5</position>
<input>
<ID>IN_0</ID>1115 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1242</ID>
<type>DA_FROM</type>
<position>386.5,6493</position>
<input>
<ID>IN_0</ID>1097 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g7</lparam></gate>
<gate>
<ID>1243</ID>
<type>AO_XNOR2</type>
<position>415.5,6496.5</position>
<input>
<ID>IN_0</ID>1113 </input>
<input>
<ID>IN_1</ID>1116 </input>
<output>
<ID>OUT</ID>1114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1244</ID>
<type>DA_FROM</type>
<position>406.5,6498.5</position>
<input>
<ID>IN_0</ID>1113 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>1245</ID>
<type>DA_FROM</type>
<position>406.5,6491</position>
<input>
<ID>IN_0</ID>1115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>1246</ID>
<type>DA_FROM</type>
<position>406.5,6494.5</position>
<input>
<ID>IN_0</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>1247</ID>
<type>DA_FROM</type>
<position>406.5,6488</position>
<input>
<ID>IN_0</ID>1117 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as7</lparam></gate>
<gate>
<ID>1248</ID>
<type>DE_TO</type>
<position>430.5,6493</position>
<input>
<ID>IN_0</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID v</lparam></gate>
<gate>
<ID>1335</ID>
<type>DA_FROM</type>
<position>226,6570</position>
<input>
<ID>IN_0</ID>856 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>1336</ID>
<type>DA_FROM</type>
<position>226,6572</position>
<input>
<ID>IN_0</ID>857 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx0</lparam></gate>
<gate>
<ID>1337</ID>
<type>DA_FROM</type>
<position>226,6574</position>
<input>
<ID>IN_0</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx0</lparam></gate>
<gate>
<ID>1338</ID>
<type>DA_FROM</type>
<position>226,6576</position>
<input>
<ID>IN_0</ID>859 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as0</lparam></gate>
<gate>
<ID>1339</ID>
<type>DA_FROM</type>
<position>226,6578</position>
<input>
<ID>IN_0</ID>863 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>1340</ID>
<type>DA_FROM</type>
<position>226,6580</position>
<input>
<ID>IN_0</ID>862 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy0</lparam></gate>
<gate>
<ID>1341</ID>
<type>DA_FROM</type>
<position>226,6582</position>
<input>
<ID>IN_0</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy0</lparam></gate>
<gate>
<ID>1342</ID>
<type>DA_FROM</type>
<position>226,6584</position>
<input>
<ID>IN_0</ID>860 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as0</lparam></gate>
<gate>
<ID>1343</ID>
<type>DE_TO</type>
<position>241.5,6577</position>
<input>
<ID>IN_0</ID>864 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa0</lparam></gate>
<gate>
<ID>1344</ID>
<type>AI_MUX_8x1</type>
<position>265.5,6577</position>
<input>
<ID>IN_0</ID>868 </input>
<input>
<ID>IN_1</ID>869 </input>
<input>
<ID>IN_2</ID>870 </input>
<input>
<ID>IN_3</ID>871 </input>
<input>
<ID>IN_4</ID>875 </input>
<input>
<ID>IN_5</ID>874 </input>
<input>
<ID>IN_6</ID>873 </input>
<input>
<ID>IN_7</ID>872 </input>
<output>
<ID>OUT</ID>876 </output>
<input>
<ID>SEL_0</ID>867 </input>
<input>
<ID>SEL_1</ID>866 </input>
<input>
<ID>SEL_2</ID>865 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1345</ID>
<type>DA_FROM</type>
<position>262.5,6586</position>
<input>
<ID>IN_0</ID>865 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1346</ID>
<type>DA_FROM</type>
<position>262.5,6588</position>
<input>
<ID>IN_0</ID>866 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1347</ID>
<type>DA_FROM</type>
<position>262.5,6590</position>
<input>
<ID>IN_0</ID>867 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1348</ID>
<type>DA_FROM</type>
<position>256.5,6570</position>
<input>
<ID>IN_0</ID>868 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>1349</ID>
<type>DA_FROM</type>
<position>256.5,6572</position>
<input>
<ID>IN_0</ID>869 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx1</lparam></gate>
<gate>
<ID>1350</ID>
<type>DA_FROM</type>
<position>256.5,6574</position>
<input>
<ID>IN_0</ID>870 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx1</lparam></gate>
<gate>
<ID>1351</ID>
<type>DA_FROM</type>
<position>256.5,6576</position>
<input>
<ID>IN_0</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as1</lparam></gate>
<gate>
<ID>1352</ID>
<type>DA_FROM</type>
<position>256.5,6578</position>
<input>
<ID>IN_0</ID>875 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>1353</ID>
<type>DA_FROM</type>
<position>256.5,6580</position>
<input>
<ID>IN_0</ID>874 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy1</lparam></gate>
<gate>
<ID>1354</ID>
<type>DA_FROM</type>
<position>256.5,6582</position>
<input>
<ID>IN_0</ID>873 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy1</lparam></gate>
<gate>
<ID>1355</ID>
<type>DA_FROM</type>
<position>256.5,6584</position>
<input>
<ID>IN_0</ID>872 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as1</lparam></gate>
<gate>
<ID>1356</ID>
<type>DE_TO</type>
<position>272.5,6577</position>
<input>
<ID>IN_0</ID>876 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa1</lparam></gate>
<gate>
<ID>1357</ID>
<type>AI_MUX_8x1</type>
<position>264.5,6553</position>
<input>
<ID>IN_0</ID>1050 </input>
<input>
<ID>IN_1</ID>1051 </input>
<input>
<ID>IN_2</ID>1052 </input>
<input>
<ID>IN_3</ID>1053 </input>
<input>
<ID>IN_4</ID>1057 </input>
<input>
<ID>IN_5</ID>1056 </input>
<input>
<ID>IN_6</ID>1055 </input>
<input>
<ID>IN_7</ID>1054 </input>
<output>
<ID>OUT</ID>1058 </output>
<input>
<ID>SEL_0</ID>1049 </input>
<input>
<ID>SEL_1</ID>1048 </input>
<input>
<ID>SEL_2</ID>1047 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1358</ID>
<type>DA_FROM</type>
<position>261.5,6562</position>
<input>
<ID>IN_0</ID>1047 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1359</ID>
<type>DA_FROM</type>
<position>261.5,6564</position>
<input>
<ID>IN_0</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1360</ID>
<type>DA_FROM</type>
<position>261.5,6566</position>
<input>
<ID>IN_0</ID>1049 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1361</ID>
<type>DA_FROM</type>
<position>255.5,6546</position>
<input>
<ID>IN_0</ID>1050 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>1362</ID>
<type>DA_FROM</type>
<position>255.5,6548</position>
<input>
<ID>IN_0</ID>1051 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx3</lparam></gate>
<gate>
<ID>1363</ID>
<type>DA_FROM</type>
<position>255.5,6550</position>
<input>
<ID>IN_0</ID>1052 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx3</lparam></gate>
<gate>
<ID>1364</ID>
<type>DA_FROM</type>
<position>255.5,6552</position>
<input>
<ID>IN_0</ID>1053 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as3</lparam></gate>
<gate>
<ID>1365</ID>
<type>DA_FROM</type>
<position>255.5,6554</position>
<input>
<ID>IN_0</ID>1057 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>1366</ID>
<type>DA_FROM</type>
<position>255.5,6556</position>
<input>
<ID>IN_0</ID>1056 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy3</lparam></gate>
<gate>
<ID>1367</ID>
<type>DA_FROM</type>
<position>255.5,6558</position>
<input>
<ID>IN_0</ID>1055 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy3</lparam></gate>
<gate>
<ID>1368</ID>
<type>DA_FROM</type>
<position>255.5,6560</position>
<input>
<ID>IN_0</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as3</lparam></gate>
<gate>
<ID>1369</ID>
<type>DE_TO</type>
<position>271.5,6553</position>
<input>
<ID>IN_0</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa3</lparam></gate>
<gate>
<ID>1370</ID>
<type>AI_MUX_8x1</type>
<position>234,6553</position>
<input>
<ID>IN_0</ID>1038 </input>
<input>
<ID>IN_1</ID>1039 </input>
<input>
<ID>IN_2</ID>1040 </input>
<input>
<ID>IN_3</ID>1041 </input>
<input>
<ID>IN_4</ID>1045 </input>
<input>
<ID>IN_5</ID>1044 </input>
<input>
<ID>IN_6</ID>1043 </input>
<input>
<ID>IN_7</ID>1042 </input>
<output>
<ID>OUT</ID>1046 </output>
<input>
<ID>SEL_0</ID>936 </input>
<input>
<ID>SEL_1</ID>931 </input>
<input>
<ID>SEL_2</ID>877 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1371</ID>
<type>DA_FROM</type>
<position>231,6562</position>
<input>
<ID>IN_0</ID>877 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1372</ID>
<type>DA_FROM</type>
<position>231,6564</position>
<input>
<ID>IN_0</ID>931 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1373</ID>
<type>DA_FROM</type>
<position>231,6566</position>
<input>
<ID>IN_0</ID>936 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1374</ID>
<type>DA_FROM</type>
<position>225,6546</position>
<input>
<ID>IN_0</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>1375</ID>
<type>DA_FROM</type>
<position>225,6548</position>
<input>
<ID>IN_0</ID>1039 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx2</lparam></gate>
<gate>
<ID>1376</ID>
<type>DA_FROM</type>
<position>225,6550</position>
<input>
<ID>IN_0</ID>1040 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx2</lparam></gate>
<gate>
<ID>1377</ID>
<type>DA_FROM</type>
<position>225,6552</position>
<input>
<ID>IN_0</ID>1041 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as2</lparam></gate>
<gate>
<ID>1378</ID>
<type>DA_FROM</type>
<position>225,6554</position>
<input>
<ID>IN_0</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>1379</ID>
<type>DA_FROM</type>
<position>225,6556</position>
<input>
<ID>IN_0</ID>1044 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy2</lparam></gate>
<gate>
<ID>1380</ID>
<type>DA_FROM</type>
<position>225,6558</position>
<input>
<ID>IN_0</ID>1043 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy2</lparam></gate>
<gate>
<ID>1381</ID>
<type>DA_FROM</type>
<position>225,6560</position>
<input>
<ID>IN_0</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as2</lparam></gate>
<gate>
<ID>1382</ID>
<type>DE_TO</type>
<position>240.5,6553</position>
<input>
<ID>IN_0</ID>1046 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa2</lparam></gate>
<gate>
<ID>1383</ID>
<type>AI_MUX_8x1</type>
<position>264.5,6528.5</position>
<input>
<ID>IN_0</ID>1074 </input>
<input>
<ID>IN_1</ID>1075 </input>
<input>
<ID>IN_2</ID>1076 </input>
<input>
<ID>IN_3</ID>1077 </input>
<input>
<ID>IN_4</ID>1081 </input>
<input>
<ID>IN_5</ID>1080 </input>
<input>
<ID>IN_6</ID>1079 </input>
<input>
<ID>IN_7</ID>1078 </input>
<output>
<ID>OUT</ID>1082 </output>
<input>
<ID>SEL_0</ID>1073 </input>
<input>
<ID>SEL_1</ID>1072 </input>
<input>
<ID>SEL_2</ID>1071 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1384</ID>
<type>DA_FROM</type>
<position>261.5,6537.5</position>
<input>
<ID>IN_0</ID>1071 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1385</ID>
<type>DA_FROM</type>
<position>261.5,6539.5</position>
<input>
<ID>IN_0</ID>1072 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1386</ID>
<type>DA_FROM</type>
<position>261.5,6541.5</position>
<input>
<ID>IN_0</ID>1073 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1387</ID>
<type>DA_FROM</type>
<position>255.5,6521.5</position>
<input>
<ID>IN_0</ID>1074 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>1388</ID>
<type>DA_FROM</type>
<position>255.5,6523.5</position>
<input>
<ID>IN_0</ID>1075 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx5</lparam></gate>
<gate>
<ID>1389</ID>
<type>DA_FROM</type>
<position>255.5,6525.5</position>
<input>
<ID>IN_0</ID>1076 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx5</lparam></gate>
<gate>
<ID>1390</ID>
<type>DA_FROM</type>
<position>255.5,6527.5</position>
<input>
<ID>IN_0</ID>1077 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as5</lparam></gate>
<gate>
<ID>1391</ID>
<type>DA_FROM</type>
<position>255.5,6529.5</position>
<input>
<ID>IN_0</ID>1081 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>1392</ID>
<type>DA_FROM</type>
<position>255.5,6531.5</position>
<input>
<ID>IN_0</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy5</lparam></gate>
<gate>
<ID>1393</ID>
<type>DA_FROM</type>
<position>255.5,6533.5</position>
<input>
<ID>IN_0</ID>1079 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy5</lparam></gate>
<gate>
<ID>1394</ID>
<type>DA_FROM</type>
<position>255.5,6535.5</position>
<input>
<ID>IN_0</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as5</lparam></gate>
<gate>
<ID>1395</ID>
<type>DE_TO</type>
<position>271.5,6528.5</position>
<input>
<ID>IN_0</ID>1082 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa5</lparam></gate>
<gate>
<ID>1396</ID>
<type>AI_MUX_8x1</type>
<position>234,6528.5</position>
<input>
<ID>IN_0</ID>1062 </input>
<input>
<ID>IN_1</ID>1063 </input>
<input>
<ID>IN_2</ID>1064 </input>
<input>
<ID>IN_3</ID>1065 </input>
<input>
<ID>IN_4</ID>1069 </input>
<input>
<ID>IN_5</ID>1068 </input>
<input>
<ID>IN_6</ID>1067 </input>
<input>
<ID>IN_7</ID>1066 </input>
<output>
<ID>OUT</ID>1070 </output>
<input>
<ID>SEL_0</ID>1061 </input>
<input>
<ID>SEL_1</ID>1060 </input>
<input>
<ID>SEL_2</ID>1059 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1397</ID>
<type>DA_FROM</type>
<position>231,6537.5</position>
<input>
<ID>IN_0</ID>1059 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1398</ID>
<type>DA_FROM</type>
<position>231,6539.5</position>
<input>
<ID>IN_0</ID>1060 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1399</ID>
<type>DA_FROM</type>
<position>231,6541.5</position>
<input>
<ID>IN_0</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1400</ID>
<type>DA_FROM</type>
<position>225,6521.5</position>
<input>
<ID>IN_0</ID>1062 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>1401</ID>
<type>DA_FROM</type>
<position>225,6523.5</position>
<input>
<ID>IN_0</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx4</lparam></gate>
<gate>
<ID>1402</ID>
<type>DA_FROM</type>
<position>225,6525.5</position>
<input>
<ID>IN_0</ID>1064 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx4</lparam></gate>
<gate>
<ID>1403</ID>
<type>DA_FROM</type>
<position>225,6527.5</position>
<input>
<ID>IN_0</ID>1065 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as4</lparam></gate>
<gate>
<ID>1404</ID>
<type>DA_FROM</type>
<position>225,6529.5</position>
<input>
<ID>IN_0</ID>1069 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>1405</ID>
<type>DA_FROM</type>
<position>225,6531.5</position>
<input>
<ID>IN_0</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy4</lparam></gate>
<gate>
<ID>1406</ID>
<type>DA_FROM</type>
<position>225,6533.5</position>
<input>
<ID>IN_0</ID>1067 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy4</lparam></gate>
<gate>
<ID>1407</ID>
<type>DA_FROM</type>
<position>225,6535.5</position>
<input>
<ID>IN_0</ID>1066 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as4</lparam></gate>
<gate>
<ID>1408</ID>
<type>DE_TO</type>
<position>240.5,6528.5</position>
<input>
<ID>IN_0</ID>1070 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa4</lparam></gate>
<gate>
<ID>1409</ID>
<type>AI_MUX_8x1</type>
<position>264.5,6504.5</position>
<input>
<ID>IN_0</ID>1135 </input>
<input>
<ID>IN_1</ID>1161 </input>
<input>
<ID>IN_2</ID>1178 </input>
<input>
<ID>IN_3</ID>1179 </input>
<input>
<ID>IN_4</ID>1183 </input>
<input>
<ID>IN_5</ID>1182 </input>
<input>
<ID>IN_6</ID>1181 </input>
<input>
<ID>IN_7</ID>1180 </input>
<output>
<ID>OUT</ID>1184 </output>
<input>
<ID>SEL_0</ID>1098 </input>
<input>
<ID>SEL_1</ID>1096 </input>
<input>
<ID>SEL_2</ID>1095 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1410</ID>
<type>DA_FROM</type>
<position>261.5,6513.5</position>
<input>
<ID>IN_0</ID>1095 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1411</ID>
<type>DA_FROM</type>
<position>261.5,6515.5</position>
<input>
<ID>IN_0</ID>1096 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1412</ID>
<type>DA_FROM</type>
<position>261.5,6517.5</position>
<input>
<ID>IN_0</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1413</ID>
<type>DA_FROM</type>
<position>255.5,6497.5</position>
<input>
<ID>IN_0</ID>1135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>1414</ID>
<type>DA_FROM</type>
<position>255.5,6499.5</position>
<input>
<ID>IN_0</ID>1161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx7</lparam></gate>
<gate>
<ID>1415</ID>
<type>DA_FROM</type>
<position>255.5,6501.5</position>
<input>
<ID>IN_0</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx7</lparam></gate>
<gate>
<ID>1416</ID>
<type>DA_FROM</type>
<position>255.5,6503.5</position>
<input>
<ID>IN_0</ID>1179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as7</lparam></gate>
<gate>
<ID>1417</ID>
<type>DA_FROM</type>
<position>255.5,6505.5</position>
<input>
<ID>IN_0</ID>1183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>1418</ID>
<type>DA_FROM</type>
<position>255.5,6507.5</position>
<input>
<ID>IN_0</ID>1182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy7</lparam></gate>
<gate>
<ID>1419</ID>
<type>DA_FROM</type>
<position>255.5,6509.5</position>
<input>
<ID>IN_0</ID>1181 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy7</lparam></gate>
<gate>
<ID>1420</ID>
<type>DA_FROM</type>
<position>255.5,6511.5</position>
<input>
<ID>IN_0</ID>1180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as7</lparam></gate>
<gate>
<ID>1421</ID>
<type>DE_TO</type>
<position>271.5,6504.5</position>
<input>
<ID>IN_0</ID>1184 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa7</lparam></gate>
<gate>
<ID>1422</ID>
<type>AI_MUX_8x1</type>
<position>234,6504.5</position>
<input>
<ID>IN_0</ID>1086 </input>
<input>
<ID>IN_1</ID>1087 </input>
<input>
<ID>IN_2</ID>1088 </input>
<input>
<ID>IN_3</ID>1089 </input>
<input>
<ID>IN_4</ID>1093 </input>
<input>
<ID>IN_5</ID>1092 </input>
<input>
<ID>IN_6</ID>1091 </input>
<input>
<ID>IN_7</ID>1090 </input>
<output>
<ID>OUT</ID>1094 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<input>
<ID>SEL_1</ID>1084 </input>
<input>
<ID>SEL_2</ID>1083 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1423</ID>
<type>DA_FROM</type>
<position>231,6513.5</position>
<input>
<ID>IN_0</ID>1083 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1424</ID>
<type>DA_FROM</type>
<position>231,6515.5</position>
<input>
<ID>IN_0</ID>1084 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1425</ID>
<type>DA_FROM</type>
<position>231,6517.5</position>
<input>
<ID>IN_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1426</ID>
<type>DA_FROM</type>
<position>225,6497.5</position>
<input>
<ID>IN_0</ID>1086 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>1427</ID>
<type>DA_FROM</type>
<position>225,6499.5</position>
<input>
<ID>IN_0</ID>1087 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incx6</lparam></gate>
<gate>
<ID>1428</ID>
<type>DA_FROM</type>
<position>225,6501.5</position>
<input>
<ID>IN_0</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decx6</lparam></gate>
<gate>
<ID>1429</ID>
<type>DA_FROM</type>
<position>225,6503.5</position>
<input>
<ID>IN_0</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as6</lparam></gate>
<gate>
<ID>1430</ID>
<type>DA_FROM</type>
<position>225,6505.5</position>
<input>
<ID>IN_0</ID>1093 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>1431</ID>
<type>DA_FROM</type>
<position>225,6507.5</position>
<input>
<ID>IN_0</ID>1092 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incy5</lparam></gate>
<gate>
<ID>1432</ID>
<type>DA_FROM</type>
<position>225,6509.5</position>
<input>
<ID>IN_0</ID>1091 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID decy5</lparam></gate>
<gate>
<ID>1433</ID>
<type>DA_FROM</type>
<position>225,6511.5</position>
<input>
<ID>IN_0</ID>1090 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID as6</lparam></gate>
<gate>
<ID>1434</ID>
<type>DE_TO</type>
<position>240.5,6504.5</position>
<input>
<ID>IN_0</ID>1094 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID oa6</lparam></gate>
<gate>
<ID>1435</ID>
<type>AA_LABEL</type>
<position>247,6597</position>
<gparam>LABEL_TEXT Mux Operacoes Aritmeticas</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>1436</ID>
<type>AI_MUX_8x1</type>
<position>235,6577</position>
<input>
<ID>IN_0</ID>856 </input>
<input>
<ID>IN_1</ID>857 </input>
<input>
<ID>IN_2</ID>858 </input>
<input>
<ID>IN_3</ID>859 </input>
<input>
<ID>IN_4</ID>863 </input>
<input>
<ID>IN_5</ID>862 </input>
<input>
<ID>IN_6</ID>861 </input>
<input>
<ID>IN_7</ID>860 </input>
<output>
<ID>OUT</ID>864 </output>
<input>
<ID>SEL_0</ID>855 </input>
<input>
<ID>SEL_1</ID>854 </input>
<input>
<ID>SEL_2</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1437</ID>
<type>DA_FROM</type>
<position>232,6586</position>
<input>
<ID>IN_0</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1438</ID>
<type>DA_FROM</type>
<position>232,6588</position>
<input>
<ID>IN_0</ID>854 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1439</ID>
<type>DA_FROM</type>
<position>232,6590</position>
<input>
<ID>IN_0</ID>855 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1440</ID>
<type>DA_FROM</type>
<position>329.5,6581</position>
<input>
<ID>IN_0</ID>1202 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx1</lparam></gate>
<gate>
<ID>1441</ID>
<type>DA_FROM</type>
<position>330.5,6583</position>
<input>
<ID>IN_0</ID>1201 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMP</lparam></gate>
<gate>
<ID>1442</ID>
<type>DA_FROM</type>
<position>329.5,6575</position>
<input>
<ID>IN_0</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor1</lparam></gate>
<gate>
<ID>1443</ID>
<type>DA_FROM</type>
<position>328,6573</position>
<input>
<ID>IN_0</ID>1206 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor1</lparam></gate>
<gate>
<ID>1444</ID>
<type>DA_FROM</type>
<position>329,6570.5</position>
<input>
<ID>IN_0</ID>1207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or1</lparam></gate>
<gate>
<ID>1445</ID>
<type>DA_FROM</type>
<position>328.5,6568</position>
<input>
<ID>IN_0</ID>1208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and1</lparam></gate>
<gate>
<ID>1446</ID>
<type>DA_FROM</type>
<position>329.5,6553</position>
<input>
<ID>IN_0</ID>1226 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx3</lparam></gate>
<gate>
<ID>1447</ID>
<type>DA_FROM</type>
<position>330.5,6555</position>
<input>
<ID>IN_0</ID>1225 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMP</lparam></gate>
<gate>
<ID>1448</ID>
<type>DA_FROM</type>
<position>329.5,6547</position>
<input>
<ID>IN_0</ID>1229 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor3</lparam></gate>
<gate>
<ID>1449</ID>
<type>DA_FROM</type>
<position>328,6545</position>
<input>
<ID>IN_0</ID>1230 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor3</lparam></gate>
<gate>
<ID>1450</ID>
<type>DA_FROM</type>
<position>329,6542.5</position>
<input>
<ID>IN_0</ID>1231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or3</lparam></gate>
<gate>
<ID>1451</ID>
<type>DA_FROM</type>
<position>328.5,6540</position>
<input>
<ID>IN_0</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and3</lparam></gate>
<gate>
<ID>1452</ID>
<type>AI_MUX_8x1</type>
<position>309,6549.5</position>
<input>
<ID>IN_0</ID>1220 </input>
<input>
<ID>IN_1</ID>1219 </input>
<input>
<ID>IN_2</ID>1218 </input>
<input>
<ID>IN_3</ID>1217 </input>
<input>
<ID>IN_4</ID>1216 </input>
<input>
<ID>IN_5</ID>1215 </input>
<input>
<ID>IN_6</ID>1214 </input>
<input>
<ID>IN_7</ID>1213 </input>
<output>
<ID>OUT</ID>1209 </output>
<input>
<ID>SEL_0</ID>1211 </input>
<input>
<ID>SEL_1</ID>1210 </input>
<input>
<ID>SEL_2</ID>1212 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1453</ID>
<type>DE_TO</type>
<position>314,6549.5</position>
<input>
<ID>IN_0</ID>1209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol2</lparam></gate>
<gate>
<ID>1454</ID>
<type>DA_FROM</type>
<position>306,6559.5</position>
<input>
<ID>IN_0</ID>1210 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1455</ID>
<type>DA_FROM</type>
<position>307,6561.5</position>
<input>
<ID>IN_0</ID>1211 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1456</ID>
<type>DA_FROM</type>
<position>304.5,6557.5</position>
<input>
<ID>IN_0</ID>1212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1457</ID>
<type>DA_FROM</type>
<position>299,6549</position>
<input>
<ID>IN_0</ID>1216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand2</lparam></gate>
<gate>
<ID>1458</ID>
<type>DA_FROM</type>
<position>298,6551</position>
<input>
<ID>IN_0</ID>1215 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor2</lparam></gate>
<gate>
<ID>1459</ID>
<type>DA_FROM</type>
<position>300,6553</position>
<input>
<ID>IN_0</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx2</lparam></gate>
<gate>
<ID>1460</ID>
<type>DA_FROM</type>
<position>301,6555</position>
<input>
<ID>IN_0</ID>1213 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMP</lparam></gate>
<gate>
<ID>1461</ID>
<type>DA_FROM</type>
<position>300,6547</position>
<input>
<ID>IN_0</ID>1217 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor2</lparam></gate>
<gate>
<ID>1462</ID>
<type>DA_FROM</type>
<position>298.5,6545</position>
<input>
<ID>IN_0</ID>1218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor2</lparam></gate>
<gate>
<ID>1463</ID>
<type>DA_FROM</type>
<position>299.5,6542.5</position>
<input>
<ID>IN_0</ID>1219 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or2</lparam></gate>
<gate>
<ID>1464</ID>
<type>DA_FROM</type>
<position>299,6540</position>
<input>
<ID>IN_0</ID>1220 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and2</lparam></gate>
<gate>
<ID>1465</ID>
<type>AI_MUX_8x1</type>
<position>338.5,6549.5</position>
<input>
<ID>IN_0</ID>1232 </input>
<input>
<ID>IN_1</ID>1231 </input>
<input>
<ID>IN_2</ID>1230 </input>
<input>
<ID>IN_3</ID>1229 </input>
<input>
<ID>IN_4</ID>1228 </input>
<input>
<ID>IN_5</ID>1227 </input>
<input>
<ID>IN_6</ID>1226 </input>
<input>
<ID>IN_7</ID>1225 </input>
<output>
<ID>OUT</ID>1221 </output>
<input>
<ID>SEL_0</ID>1223 </input>
<input>
<ID>SEL_1</ID>1222 </input>
<input>
<ID>SEL_2</ID>1224 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1466</ID>
<type>DE_TO</type>
<position>343.5,6549.5</position>
<input>
<ID>IN_0</ID>1221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol3</lparam></gate>
<gate>
<ID>1467</ID>
<type>DA_FROM</type>
<position>335.5,6559.5</position>
<input>
<ID>IN_0</ID>1222 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1468</ID>
<type>DA_FROM</type>
<position>336.5,6561.5</position>
<input>
<ID>IN_0</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1469</ID>
<type>DA_FROM</type>
<position>334,6557.5</position>
<input>
<ID>IN_0</ID>1224 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1470</ID>
<type>DA_FROM</type>
<position>328.5,6549</position>
<input>
<ID>IN_0</ID>1228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand3</lparam></gate>
<gate>
<ID>1471</ID>
<type>DA_FROM</type>
<position>327.5,6551</position>
<input>
<ID>IN_0</ID>1227 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor3</lparam></gate>
<gate>
<ID>1472</ID>
<type>DA_FROM</type>
<position>329.5,6525</position>
<input>
<ID>IN_0</ID>1250 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx5</lparam></gate>
<gate>
<ID>1473</ID>
<type>DA_FROM</type>
<position>330.5,6527</position>
<input>
<ID>IN_0</ID>1249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMP</lparam></gate>
<gate>
<ID>1474</ID>
<type>DA_FROM</type>
<position>329.5,6519</position>
<input>
<ID>IN_0</ID>1253 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor5</lparam></gate>
<gate>
<ID>1475</ID>
<type>DA_FROM</type>
<position>328,6517</position>
<input>
<ID>IN_0</ID>1254 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor5</lparam></gate>
<gate>
<ID>1476</ID>
<type>DA_FROM</type>
<position>329,6514.5</position>
<input>
<ID>IN_0</ID>1255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or5</lparam></gate>
<gate>
<ID>1477</ID>
<type>DA_FROM</type>
<position>328.5,6512</position>
<input>
<ID>IN_0</ID>1256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and5</lparam></gate>
<gate>
<ID>1478</ID>
<type>DA_FROM</type>
<position>329.5,6497</position>
<input>
<ID>IN_0</ID>1274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx7</lparam></gate>
<gate>
<ID>1479</ID>
<type>DA_FROM</type>
<position>330.5,6499</position>
<input>
<ID>IN_0</ID>1273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMP</lparam></gate>
<gate>
<ID>1480</ID>
<type>DA_FROM</type>
<position>329.5,6491</position>
<input>
<ID>IN_0</ID>1277 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor7</lparam></gate>
<gate>
<ID>1481</ID>
<type>DA_FROM</type>
<position>328,6489</position>
<input>
<ID>IN_0</ID>1278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor7</lparam></gate>
<gate>
<ID>1482</ID>
<type>DA_FROM</type>
<position>329,6486.5</position>
<input>
<ID>IN_0</ID>1279 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or7</lparam></gate>
<gate>
<ID>1483</ID>
<type>DA_FROM</type>
<position>328.5,6484</position>
<input>
<ID>IN_0</ID>1280 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and7</lparam></gate>
<gate>
<ID>1484</ID>
<type>AI_MUX_8x1</type>
<position>309,6493.5</position>
<input>
<ID>IN_0</ID>1268 </input>
<input>
<ID>IN_1</ID>1267 </input>
<input>
<ID>IN_2</ID>1266 </input>
<input>
<ID>IN_3</ID>1265 </input>
<input>
<ID>IN_4</ID>1264 </input>
<input>
<ID>IN_5</ID>1263 </input>
<input>
<ID>IN_6</ID>1262 </input>
<input>
<ID>IN_7</ID>1261 </input>
<output>
<ID>OUT</ID>1257 </output>
<input>
<ID>SEL_0</ID>1259 </input>
<input>
<ID>SEL_1</ID>1258 </input>
<input>
<ID>SEL_2</ID>1260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1485</ID>
<type>DE_TO</type>
<position>314,6493.5</position>
<input>
<ID>IN_0</ID>1257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol6</lparam></gate>
<gate>
<ID>1486</ID>
<type>DA_FROM</type>
<position>306,6503.5</position>
<input>
<ID>IN_0</ID>1258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1487</ID>
<type>DA_FROM</type>
<position>307,6505.5</position>
<input>
<ID>IN_0</ID>1259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1488</ID>
<type>DA_FROM</type>
<position>304.5,6501.5</position>
<input>
<ID>IN_0</ID>1260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1489</ID>
<type>DA_FROM</type>
<position>299,6493</position>
<input>
<ID>IN_0</ID>1264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand6</lparam></gate>
<gate>
<ID>1490</ID>
<type>DA_FROM</type>
<position>298,6495</position>
<input>
<ID>IN_0</ID>1263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor6</lparam></gate>
<gate>
<ID>1491</ID>
<type>DA_FROM</type>
<position>300,6497</position>
<input>
<ID>IN_0</ID>1262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx6</lparam></gate>
<gate>
<ID>1492</ID>
<type>DA_FROM</type>
<position>301,6499</position>
<input>
<ID>IN_0</ID>1261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMP</lparam></gate>
<gate>
<ID>1493</ID>
<type>DA_FROM</type>
<position>300,6491</position>
<input>
<ID>IN_0</ID>1265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor6</lparam></gate>
<gate>
<ID>1494</ID>
<type>DA_FROM</type>
<position>298.5,6489</position>
<input>
<ID>IN_0</ID>1266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor6</lparam></gate>
<gate>
<ID>1495</ID>
<type>DA_FROM</type>
<position>299.5,6486.5</position>
<input>
<ID>IN_0</ID>1267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or6</lparam></gate>
<gate>
<ID>1496</ID>
<type>DA_FROM</type>
<position>299,6484</position>
<input>
<ID>IN_0</ID>1268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and6</lparam></gate>
<gate>
<ID>1497</ID>
<type>AI_MUX_8x1</type>
<position>338.5,6493.5</position>
<input>
<ID>IN_0</ID>1280 </input>
<input>
<ID>IN_1</ID>1279 </input>
<input>
<ID>IN_2</ID>1278 </input>
<input>
<ID>IN_3</ID>1277 </input>
<input>
<ID>IN_4</ID>1276 </input>
<input>
<ID>IN_5</ID>1275 </input>
<input>
<ID>IN_6</ID>1274 </input>
<input>
<ID>IN_7</ID>1273 </input>
<output>
<ID>OUT</ID>1269 </output>
<input>
<ID>SEL_0</ID>1271 </input>
<input>
<ID>SEL_1</ID>1270 </input>
<input>
<ID>SEL_2</ID>1272 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1498</ID>
<type>DE_TO</type>
<position>343.5,6493.5</position>
<input>
<ID>IN_0</ID>1269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol7</lparam></gate>
<gate>
<ID>1499</ID>
<type>DA_FROM</type>
<position>335.5,6503.5</position>
<input>
<ID>IN_0</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1500</ID>
<type>DA_FROM</type>
<position>336.5,6505.5</position>
<input>
<ID>IN_0</ID>1271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1501</ID>
<type>DA_FROM</type>
<position>334,6501.5</position>
<input>
<ID>IN_0</ID>1272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1502</ID>
<type>DA_FROM</type>
<position>328.5,6493</position>
<input>
<ID>IN_0</ID>1276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand7</lparam></gate>
<gate>
<ID>1503</ID>
<type>DA_FROM</type>
<position>327.5,6495</position>
<input>
<ID>IN_0</ID>1275 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor7</lparam></gate>
<gate>
<ID>1504</ID>
<type>AI_MUX_8x1</type>
<position>309,6521.5</position>
<input>
<ID>IN_0</ID>1244 </input>
<input>
<ID>IN_1</ID>1243 </input>
<input>
<ID>IN_2</ID>1242 </input>
<input>
<ID>IN_3</ID>1241 </input>
<input>
<ID>IN_4</ID>1240 </input>
<input>
<ID>IN_5</ID>1239 </input>
<input>
<ID>IN_6</ID>1238 </input>
<input>
<ID>IN_7</ID>1237 </input>
<output>
<ID>OUT</ID>1233 </output>
<input>
<ID>SEL_0</ID>1235 </input>
<input>
<ID>SEL_1</ID>1234 </input>
<input>
<ID>SEL_2</ID>1236 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1505</ID>
<type>DE_TO</type>
<position>314,6521.5</position>
<input>
<ID>IN_0</ID>1233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol4</lparam></gate>
<gate>
<ID>1506</ID>
<type>DA_FROM</type>
<position>306,6531.5</position>
<input>
<ID>IN_0</ID>1234 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1507</ID>
<type>DA_FROM</type>
<position>307,6533.5</position>
<input>
<ID>IN_0</ID>1235 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1508</ID>
<type>DA_FROM</type>
<position>304.5,6529.5</position>
<input>
<ID>IN_0</ID>1236 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1509</ID>
<type>DA_FROM</type>
<position>299,6521</position>
<input>
<ID>IN_0</ID>1240 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand4</lparam></gate>
<gate>
<ID>1510</ID>
<type>DA_FROM</type>
<position>298,6523</position>
<input>
<ID>IN_0</ID>1239 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor4</lparam></gate>
<gate>
<ID>1511</ID>
<type>DA_FROM</type>
<position>300,6525</position>
<input>
<ID>IN_0</ID>1238 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx4</lparam></gate>
<gate>
<ID>1512</ID>
<type>DA_FROM</type>
<position>301,6527</position>
<input>
<ID>IN_0</ID>1237 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMP</lparam></gate>
<gate>
<ID>1513</ID>
<type>DA_FROM</type>
<position>300,6519</position>
<input>
<ID>IN_0</ID>1241 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor4</lparam></gate>
<gate>
<ID>1514</ID>
<type>DA_FROM</type>
<position>298.5,6517</position>
<input>
<ID>IN_0</ID>1242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor4</lparam></gate>
<gate>
<ID>1515</ID>
<type>DA_FROM</type>
<position>299.5,6514.5</position>
<input>
<ID>IN_0</ID>1243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or4</lparam></gate>
<gate>
<ID>1516</ID>
<type>DA_FROM</type>
<position>299,6512</position>
<input>
<ID>IN_0</ID>1244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and4</lparam></gate>
<gate>
<ID>1517</ID>
<type>AI_MUX_8x1</type>
<position>338.5,6521.5</position>
<input>
<ID>IN_0</ID>1256 </input>
<input>
<ID>IN_1</ID>1255 </input>
<input>
<ID>IN_2</ID>1254 </input>
<input>
<ID>IN_3</ID>1253 </input>
<input>
<ID>IN_4</ID>1252 </input>
<input>
<ID>IN_5</ID>1251 </input>
<input>
<ID>IN_6</ID>1250 </input>
<input>
<ID>IN_7</ID>1249 </input>
<output>
<ID>OUT</ID>1245 </output>
<input>
<ID>SEL_0</ID>1247 </input>
<input>
<ID>SEL_1</ID>1246 </input>
<input>
<ID>SEL_2</ID>1248 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1518</ID>
<type>DE_TO</type>
<position>343.5,6521.5</position>
<input>
<ID>IN_0</ID>1245 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol5</lparam></gate>
<gate>
<ID>1519</ID>
<type>DA_FROM</type>
<position>335.5,6531.5</position>
<input>
<ID>IN_0</ID>1246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1520</ID>
<type>DA_FROM</type>
<position>336.5,6533.5</position>
<input>
<ID>IN_0</ID>1247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1521</ID>
<type>DA_FROM</type>
<position>334,6529.5</position>
<input>
<ID>IN_0</ID>1248 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1522</ID>
<type>DA_FROM</type>
<position>328.5,6521</position>
<input>
<ID>IN_0</ID>1252 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand5</lparam></gate>
<gate>
<ID>1523</ID>
<type>DA_FROM</type>
<position>327.5,6523</position>
<input>
<ID>IN_0</ID>1251 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor5</lparam></gate>
<gate>
<ID>1524</ID>
<type>AA_LABEL</type>
<position>321,6597.5</position>
<gparam>LABEL_TEXT Mux Operacoes Logicas</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1525</ID>
<type>AI_MUX_8x1</type>
<position>309,6577.5</position>
<input>
<ID>IN_0</ID>1196 </input>
<input>
<ID>IN_1</ID>1195 </input>
<input>
<ID>IN_2</ID>1194 </input>
<input>
<ID>IN_3</ID>1193 </input>
<input>
<ID>IN_4</ID>1192 </input>
<input>
<ID>IN_5</ID>1191 </input>
<input>
<ID>IN_6</ID>1190 </input>
<input>
<ID>IN_7</ID>1189 </input>
<output>
<ID>OUT</ID>1185 </output>
<input>
<ID>SEL_0</ID>1187 </input>
<input>
<ID>SEL_1</ID>1186 </input>
<input>
<ID>SEL_2</ID>1188 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1526</ID>
<type>DE_TO</type>
<position>314,6577.5</position>
<input>
<ID>IN_0</ID>1185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol0</lparam></gate>
<gate>
<ID>1527</ID>
<type>DA_FROM</type>
<position>306,6587.5</position>
<input>
<ID>IN_0</ID>1186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1528</ID>
<type>DA_FROM</type>
<position>307,6589.5</position>
<input>
<ID>IN_0</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1529</ID>
<type>DA_FROM</type>
<position>304.5,6585.5</position>
<input>
<ID>IN_0</ID>1188 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1530</ID>
<type>DA_FROM</type>
<position>299,6577</position>
<input>
<ID>IN_0</ID>1192 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand0</lparam></gate>
<gate>
<ID>1531</ID>
<type>DA_FROM</type>
<position>298,6579</position>
<input>
<ID>IN_0</ID>1191 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor0</lparam></gate>
<gate>
<ID>1532</ID>
<type>DA_FROM</type>
<position>300,6581</position>
<input>
<ID>IN_0</ID>1190 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID notx0</lparam></gate>
<gate>
<ID>1533</ID>
<type>DA_FROM</type>
<position>301,6583</position>
<input>
<ID>IN_0</ID>1189 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMP</lparam></gate>
<gate>
<ID>1534</ID>
<type>DA_FROM</type>
<position>300,6575</position>
<input>
<ID>IN_0</ID>1193 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xnor0</lparam></gate>
<gate>
<ID>1535</ID>
<type>DA_FROM</type>
<position>298.5,6573</position>
<input>
<ID>IN_0</ID>1194 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID xor0</lparam></gate>
<gate>
<ID>1536</ID>
<type>DA_FROM</type>
<position>299.5,6570.5</position>
<input>
<ID>IN_0</ID>1195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID or0</lparam></gate>
<gate>
<ID>1537</ID>
<type>DA_FROM</type>
<position>299,6568</position>
<input>
<ID>IN_0</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID and0</lparam></gate>
<gate>
<ID>1538</ID>
<type>AI_MUX_8x1</type>
<position>338.5,6577.5</position>
<input>
<ID>IN_0</ID>1208 </input>
<input>
<ID>IN_1</ID>1207 </input>
<input>
<ID>IN_2</ID>1206 </input>
<input>
<ID>IN_3</ID>1205 </input>
<input>
<ID>IN_4</ID>1204 </input>
<input>
<ID>IN_5</ID>1203 </input>
<input>
<ID>IN_6</ID>1202 </input>
<input>
<ID>IN_7</ID>1201 </input>
<output>
<ID>OUT</ID>1197 </output>
<input>
<ID>SEL_0</ID>1199 </input>
<input>
<ID>SEL_1</ID>1198 </input>
<input>
<ID>SEL_2</ID>1200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1539</ID>
<type>DE_TO</type>
<position>343.5,6577.5</position>
<input>
<ID>IN_0</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ol1</lparam></gate>
<gate>
<ID>1540</ID>
<type>DA_FROM</type>
<position>335.5,6587.5</position>
<input>
<ID>IN_0</ID>1198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>1541</ID>
<type>DA_FROM</type>
<position>336.5,6589.5</position>
<input>
<ID>IN_0</ID>1199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>1542</ID>
<type>DA_FROM</type>
<position>334,6585.5</position>
<input>
<ID>IN_0</ID>1200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s2</lparam></gate>
<gate>
<ID>1543</ID>
<type>DA_FROM</type>
<position>328.5,6577</position>
<input>
<ID>IN_0</ID>1204 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nand0</lparam></gate>
<gate>
<ID>1544</ID>
<type>DA_FROM</type>
<position>327.5,6579</position>
<input>
<ID>IN_0</ID>1203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nor1</lparam></gate>
<gate>
<ID>1546</ID>
<type>AA_LABEL</type>
<position>264.5,6611</position>
<gparam>LABEL_TEXT MULTIPLEXADORES</gparam>
<gparam>TEXT_HEIGHT 7</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1547</ID>
<type>DE_TO</type>
<position>403.5,6579.5</position>
<input>
<ID>IN_0</ID>1298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g7</lparam></gate>
<gate>
<ID>1548</ID>
<type>DE_TO</type>
<position>403.5,6574.5</position>
<input>
<ID>IN_0</ID>1299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g6</lparam></gate>
<gate>
<ID>1549</ID>
<type>DE_TO</type>
<position>403.5,6569.5</position>
<input>
<ID>IN_0</ID>1300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g5</lparam></gate>
<gate>
<ID>1550</ID>
<type>DE_TO</type>
<position>403.5,6564.5</position>
<input>
<ID>IN_0</ID>1301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g4</lparam></gate>
<gate>
<ID>1551</ID>
<type>DE_TO</type>
<position>403.5,6559.5</position>
<input>
<ID>IN_0</ID>1302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g3</lparam></gate>
<gate>
<ID>1552</ID>
<type>DE_TO</type>
<position>403,6554.5</position>
<input>
<ID>IN_0</ID>1303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g2</lparam></gate>
<gate>
<ID>1553</ID>
<type>DE_TO</type>
<position>403,6549.5</position>
<input>
<ID>IN_0</ID>1304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g1</lparam></gate>
<gate>
<ID>1554</ID>
<type>DE_TO</type>
<position>403,6544.5</position>
<input>
<ID>IN_0</ID>1305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g0</lparam></gate>
<gate>
<ID>1555</ID>
<type>AA_MUX_2x1</type>
<position>393.5,6579.5</position>
<input>
<ID>IN_0</ID>1281 </input>
<input>
<ID>IN_1</ID>1297 </input>
<output>
<ID>OUT</ID>1298 </output>
<input>
<ID>SEL_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,6501.5,259.5,6503</points>
<intersection>6501.5 2</intersection>
<intersection>6503 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,6503,261.5,6503</points>
<connection>
<GID>1409</GID>
<name>IN_2</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,6501.5,259.5,6501.5</points>
<connection>
<GID>1415</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>257.5,6503.5,259.5,6503.5</points>
<connection>
<GID>1416</GID>
<name>IN_0</name></connection>
<intersection>259.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>259.5,6503.5,259.5,6504</points>
<intersection>6503.5 1</intersection>
<intersection>6504 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,6504,261.5,6504</points>
<connection>
<GID>1409</GID>
<name>IN_3</name></connection>
<intersection>259.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,6508,260.5,6511.5</points>
<intersection>6508 1</intersection>
<intersection>6511.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,6508,261.5,6508</points>
<connection>
<GID>1409</GID>
<name>IN_7</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,6511.5,260.5,6511.5</points>
<connection>
<GID>1420</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,6507,260,6509.5</points>
<intersection>6507 1</intersection>
<intersection>6509.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,6507,261.5,6507</points>
<connection>
<GID>1409</GID>
<name>IN_6</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>257.5,6509.5,260,6509.5</points>
<connection>
<GID>1419</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>1182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,6506,259.5,6507.5</points>
<intersection>6506 2</intersection>
<intersection>6507.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,6507.5,259.5,6507.5</points>
<connection>
<GID>1418</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,6506,261.5,6506</points>
<connection>
<GID>1409</GID>
<name>IN_5</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>257.5,6505.5,259.5,6505.5</points>
<connection>
<GID>1417</GID>
<name>IN_0</name></connection>
<intersection>259.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>259.5,6505,259.5,6505.5</points>
<intersection>6505 4</intersection>
<intersection>6505.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,6505,261.5,6505</points>
<connection>
<GID>1409</GID>
<name>IN_4</name></connection>
<intersection>259.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1184</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>267.5,6504.5,269.5,6504.5</points>
<connection>
<GID>1409</GID>
<name>OUT</name></connection>
<connection>
<GID>1421</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,6577.5,312,6577.5</points>
<connection>
<GID>1525</GID>
<name>OUT</name></connection>
<connection>
<GID>1526</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,6583,309,6587.5</points>
<connection>
<GID>1525</GID>
<name>SEL_1</name></connection>
<intersection>6587.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>308,6587.5,309,6587.5</points>
<connection>
<GID>1527</GID>
<name>IN_0</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>1187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,6583,310,6589.5</points>
<connection>
<GID>1525</GID>
<name>SEL_0</name></connection>
<intersection>6589.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,6589.5,310,6589.5</points>
<connection>
<GID>1528</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>1188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,6583,308,6585.5</points>
<connection>
<GID>1525</GID>
<name>SEL_2</name></connection>
<intersection>6585.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>306.5,6585.5,308,6585.5</points>
<connection>
<GID>1529</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>1189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305.5,6581,306,6581</points>
<connection>
<GID>1525</GID>
<name>IN_7</name></connection>
<intersection>305.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>305.5,6581,305.5,6583</points>
<intersection>6581 1</intersection>
<intersection>6583 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>303,6583,305.5,6583</points>
<connection>
<GID>1533</GID>
<name>IN_0</name></connection>
<intersection>305.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>302,6580,306,6580</points>
<connection>
<GID>1525</GID>
<name>IN_6</name></connection>
<intersection>302 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>302,6580,302,6581</points>
<connection>
<GID>1532</GID>
<name>IN_0</name></connection>
<intersection>6580 1</intersection></vsegment></shape></wire>
<wire>
<ID>1191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>300,6579,306,6579</points>
<connection>
<GID>1531</GID>
<name>IN_0</name></connection>
<connection>
<GID>1525</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>300.5,6577,300.5,6577.5</points>
<intersection>6577 8</intersection>
<intersection>6577.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>300.5,6577.5,306,6577.5</points>
<intersection>300.5 0</intersection>
<intersection>306 9</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>300.5,6577,301,6577</points>
<connection>
<GID>1530</GID>
<name>IN_0</name></connection>
<intersection>300.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>306,6577.5,306,6578</points>
<connection>
<GID>1525</GID>
<name>IN_4</name></connection>
<intersection>6577.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,6575,302.5,6577</points>
<intersection>6575 4</intersection>
<intersection>6577 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,6577,306,6577</points>
<connection>
<GID>1525</GID>
<name>IN_3</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>302,6575,302.5,6575</points>
<connection>
<GID>1534</GID>
<name>IN_0</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,6573,303.5,6576</points>
<intersection>6573 2</intersection>
<intersection>6576 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,6576,306,6576</points>
<connection>
<GID>1525</GID>
<name>IN_2</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,6573,303.5,6573</points>
<connection>
<GID>1535</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,6570.5,304,6575</points>
<intersection>6570.5 2</intersection>
<intersection>6575 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,6575,306,6575</points>
<connection>
<GID>1525</GID>
<name>IN_1</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,6570.5,304,6570.5</points>
<connection>
<GID>1536</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>1196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,6568,304.5,6574</points>
<intersection>6568 2</intersection>
<intersection>6574 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,6574,306,6574</points>
<connection>
<GID>1525</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,6568,304.5,6568</points>
<connection>
<GID>1537</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,6577.5,341.5,6577.5</points>
<connection>
<GID>1538</GID>
<name>OUT</name></connection>
<connection>
<GID>1539</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338.5,6583,338.5,6587.5</points>
<connection>
<GID>1538</GID>
<name>SEL_1</name></connection>
<intersection>6587.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>337.5,6587.5,338.5,6587.5</points>
<connection>
<GID>1540</GID>
<name>IN_0</name></connection>
<intersection>338.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,6583,339.5,6589.5</points>
<connection>
<GID>1538</GID>
<name>SEL_0</name></connection>
<intersection>6589.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>338.5,6589.5,339.5,6589.5</points>
<connection>
<GID>1541</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,6583,337.5,6585.5</points>
<connection>
<GID>1538</GID>
<name>SEL_2</name></connection>
<intersection>6585.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336,6585.5,337.5,6585.5</points>
<connection>
<GID>1542</GID>
<name>IN_0</name></connection>
<intersection>337.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>335,6581,335.5,6581</points>
<connection>
<GID>1538</GID>
<name>IN_7</name></connection>
<intersection>335 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>335,6581,335,6583</points>
<intersection>6581 1</intersection>
<intersection>6583 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>332.5,6583,335,6583</points>
<connection>
<GID>1441</GID>
<name>IN_0</name></connection>
<intersection>335 3</intersection></hsegment></shape></wire>
<wire>
<ID>1202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>331.5,6580,335.5,6580</points>
<connection>
<GID>1538</GID>
<name>IN_6</name></connection>
<intersection>331.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>331.5,6580,331.5,6581</points>
<connection>
<GID>1440</GID>
<name>IN_0</name></connection>
<intersection>6580 1</intersection></vsegment></shape></wire>
<wire>
<ID>1203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329.5,6579,335.5,6579</points>
<connection>
<GID>1544</GID>
<name>IN_0</name></connection>
<connection>
<GID>1538</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,6577,330,6577.5</points>
<intersection>6577 8</intersection>
<intersection>6577.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>330,6577.5,335.5,6577.5</points>
<intersection>330 0</intersection>
<intersection>335.5 9</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>330,6577,330.5,6577</points>
<connection>
<GID>1543</GID>
<name>IN_0</name></connection>
<intersection>330 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>335.5,6577.5,335.5,6578</points>
<connection>
<GID>1538</GID>
<name>IN_4</name></connection>
<intersection>6577.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,6575,332,6577</points>
<intersection>6575 2</intersection>
<intersection>6577 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332,6577,335.5,6577</points>
<connection>
<GID>1538</GID>
<name>IN_3</name></connection>
<intersection>332 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>331.5,6575,332,6575</points>
<connection>
<GID>1442</GID>
<name>IN_0</name></connection>
<intersection>332 0</intersection></hsegment></shape></wire>
<wire>
<ID>1206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,6573,333,6576</points>
<intersection>6573 2</intersection>
<intersection>6576 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,6576,335.5,6576</points>
<connection>
<GID>1538</GID>
<name>IN_2</name></connection>
<intersection>333 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330,6573,333,6573</points>
<connection>
<GID>1443</GID>
<name>IN_0</name></connection>
<intersection>333 0</intersection></hsegment></shape></wire>
<wire>
<ID>1207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,6570.5,333.5,6575</points>
<intersection>6570.5 2</intersection>
<intersection>6575 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333.5,6575,335.5,6575</points>
<connection>
<GID>1538</GID>
<name>IN_1</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>331,6570.5,333.5,6570.5</points>
<connection>
<GID>1444</GID>
<name>IN_0</name></connection>
<intersection>333.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,6568,334,6574</points>
<intersection>6568 2</intersection>
<intersection>6574 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334,6574,335.5,6574</points>
<connection>
<GID>1538</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330.5,6568,334,6568</points>
<connection>
<GID>1445</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>1209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,6549.5,312,6549.5</points>
<connection>
<GID>1452</GID>
<name>OUT</name></connection>
<connection>
<GID>1453</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,6555,309,6559.5</points>
<connection>
<GID>1452</GID>
<name>SEL_1</name></connection>
<intersection>6559.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>308,6559.5,309,6559.5</points>
<connection>
<GID>1454</GID>
<name>IN_0</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>1211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,6555,310,6561.5</points>
<connection>
<GID>1452</GID>
<name>SEL_0</name></connection>
<intersection>6561.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,6561.5,310,6561.5</points>
<connection>
<GID>1455</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>1212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,6555,308,6557.5</points>
<connection>
<GID>1452</GID>
<name>SEL_2</name></connection>
<intersection>6557.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>306.5,6557.5,308,6557.5</points>
<connection>
<GID>1456</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>1213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305.5,6553,306,6553</points>
<connection>
<GID>1452</GID>
<name>IN_7</name></connection>
<intersection>305.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>305.5,6553,305.5,6555</points>
<intersection>6553 1</intersection>
<intersection>6555 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>303,6555,305.5,6555</points>
<connection>
<GID>1460</GID>
<name>IN_0</name></connection>
<intersection>305.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>302,6552,306,6552</points>
<connection>
<GID>1452</GID>
<name>IN_6</name></connection>
<intersection>302 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>302,6552,302,6553</points>
<connection>
<GID>1459</GID>
<name>IN_0</name></connection>
<intersection>6552 1</intersection></vsegment></shape></wire>
<wire>
<ID>1215</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>300,6551,306,6551</points>
<connection>
<GID>1458</GID>
<name>IN_0</name></connection>
<connection>
<GID>1452</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>300.5,6549,300.5,6549.5</points>
<intersection>6549 8</intersection>
<intersection>6549.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>300.5,6549.5,306,6549.5</points>
<intersection>300.5 0</intersection>
<intersection>306 9</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>300.5,6549,301,6549</points>
<connection>
<GID>1457</GID>
<name>IN_0</name></connection>
<intersection>300.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>306,6549.5,306,6550</points>
<connection>
<GID>1452</GID>
<name>IN_4</name></connection>
<intersection>6549.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,6547,302.5,6549</points>
<intersection>6547 4</intersection>
<intersection>6549 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,6549,306,6549</points>
<connection>
<GID>1452</GID>
<name>IN_3</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>302,6547,302.5,6547</points>
<connection>
<GID>1461</GID>
<name>IN_0</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,6545,303.5,6548</points>
<intersection>6545 2</intersection>
<intersection>6548 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,6548,306,6548</points>
<connection>
<GID>1452</GID>
<name>IN_2</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,6545,303.5,6545</points>
<connection>
<GID>1462</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,6542.5,304,6547</points>
<intersection>6542.5 2</intersection>
<intersection>6547 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,6547,306,6547</points>
<connection>
<GID>1452</GID>
<name>IN_1</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,6542.5,304,6542.5</points>
<connection>
<GID>1463</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>1220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,6540,304.5,6546</points>
<intersection>6540 2</intersection>
<intersection>6546 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,6546,306,6546</points>
<connection>
<GID>1452</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,6540,304.5,6540</points>
<connection>
<GID>1464</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,6549.5,341.5,6549.5</points>
<connection>
<GID>1465</GID>
<name>OUT</name></connection>
<connection>
<GID>1466</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338.5,6555,338.5,6559.5</points>
<connection>
<GID>1465</GID>
<name>SEL_1</name></connection>
<intersection>6559.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>337.5,6559.5,338.5,6559.5</points>
<connection>
<GID>1467</GID>
<name>IN_0</name></connection>
<intersection>338.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,6555,339.5,6561.5</points>
<connection>
<GID>1465</GID>
<name>SEL_0</name></connection>
<intersection>6561.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>338.5,6561.5,339.5,6561.5</points>
<connection>
<GID>1468</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,6555,337.5,6557.5</points>
<connection>
<GID>1465</GID>
<name>SEL_2</name></connection>
<intersection>6557.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336,6557.5,337.5,6557.5</points>
<connection>
<GID>1469</GID>
<name>IN_0</name></connection>
<intersection>337.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>335,6553,335.5,6553</points>
<connection>
<GID>1465</GID>
<name>IN_7</name></connection>
<intersection>335 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>335,6553,335,6555</points>
<intersection>6553 1</intersection>
<intersection>6555 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>332.5,6555,335,6555</points>
<connection>
<GID>1447</GID>
<name>IN_0</name></connection>
<intersection>335 3</intersection></hsegment></shape></wire>
<wire>
<ID>1226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>331.5,6552,335.5,6552</points>
<connection>
<GID>1465</GID>
<name>IN_6</name></connection>
<intersection>331.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>331.5,6552,331.5,6553</points>
<connection>
<GID>1446</GID>
<name>IN_0</name></connection>
<intersection>6552 1</intersection></vsegment></shape></wire>
<wire>
<ID>1227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329.5,6551,335.5,6551</points>
<connection>
<GID>1471</GID>
<name>IN_0</name></connection>
<connection>
<GID>1465</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,6549,330,6549.5</points>
<intersection>6549 8</intersection>
<intersection>6549.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>330,6549.5,335.5,6549.5</points>
<intersection>330 0</intersection>
<intersection>335.5 9</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>330,6549,330.5,6549</points>
<connection>
<GID>1470</GID>
<name>IN_0</name></connection>
<intersection>330 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>335.5,6549.5,335.5,6550</points>
<connection>
<GID>1465</GID>
<name>IN_4</name></connection>
<intersection>6549.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,6547,332,6549</points>
<intersection>6547 2</intersection>
<intersection>6549 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332,6549,335.5,6549</points>
<connection>
<GID>1465</GID>
<name>IN_3</name></connection>
<intersection>332 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>331.5,6547,332,6547</points>
<connection>
<GID>1448</GID>
<name>IN_0</name></connection>
<intersection>332 0</intersection></hsegment></shape></wire>
<wire>
<ID>1230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,6545,333,6548</points>
<intersection>6545 2</intersection>
<intersection>6548 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,6548,335.5,6548</points>
<connection>
<GID>1465</GID>
<name>IN_2</name></connection>
<intersection>333 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330,6545,333,6545</points>
<connection>
<GID>1449</GID>
<name>IN_0</name></connection>
<intersection>333 0</intersection></hsegment></shape></wire>
<wire>
<ID>1231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,6542.5,333.5,6547</points>
<intersection>6542.5 2</intersection>
<intersection>6547 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333.5,6547,335.5,6547</points>
<connection>
<GID>1465</GID>
<name>IN_1</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>331,6542.5,333.5,6542.5</points>
<connection>
<GID>1450</GID>
<name>IN_0</name></connection>
<intersection>333.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,6540,334,6546</points>
<intersection>6540 2</intersection>
<intersection>6546 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334,6546,335.5,6546</points>
<connection>
<GID>1465</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330.5,6540,334,6540</points>
<connection>
<GID>1451</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>1233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,6521.5,312,6521.5</points>
<connection>
<GID>1504</GID>
<name>OUT</name></connection>
<connection>
<GID>1505</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,6527,309,6531.5</points>
<connection>
<GID>1504</GID>
<name>SEL_1</name></connection>
<intersection>6531.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>308,6531.5,309,6531.5</points>
<connection>
<GID>1506</GID>
<name>IN_0</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>1235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,6527,310,6533.5</points>
<connection>
<GID>1504</GID>
<name>SEL_0</name></connection>
<intersection>6533.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,6533.5,310,6533.5</points>
<connection>
<GID>1507</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>1236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,6527,308,6529.5</points>
<connection>
<GID>1504</GID>
<name>SEL_2</name></connection>
<intersection>6529.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>306.5,6529.5,308,6529.5</points>
<connection>
<GID>1508</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>1237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305.5,6525,306,6525</points>
<connection>
<GID>1504</GID>
<name>IN_7</name></connection>
<intersection>305.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>305.5,6525,305.5,6527</points>
<intersection>6525 1</intersection>
<intersection>6527 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>303,6527,305.5,6527</points>
<connection>
<GID>1512</GID>
<name>IN_0</name></connection>
<intersection>305.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>302,6524,306,6524</points>
<connection>
<GID>1504</GID>
<name>IN_6</name></connection>
<intersection>302 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>302,6524,302,6525</points>
<connection>
<GID>1511</GID>
<name>IN_0</name></connection>
<intersection>6524 1</intersection></vsegment></shape></wire>
<wire>
<ID>1239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>300,6523,306,6523</points>
<connection>
<GID>1510</GID>
<name>IN_0</name></connection>
<connection>
<GID>1504</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>300.5,6521,300.5,6521.5</points>
<intersection>6521 8</intersection>
<intersection>6521.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>300.5,6521.5,306,6521.5</points>
<intersection>300.5 0</intersection>
<intersection>306 9</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>300.5,6521,301,6521</points>
<connection>
<GID>1509</GID>
<name>IN_0</name></connection>
<intersection>300.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>306,6521.5,306,6522</points>
<connection>
<GID>1504</GID>
<name>IN_4</name></connection>
<intersection>6521.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,6519,302.5,6521</points>
<intersection>6519 4</intersection>
<intersection>6521 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,6521,306,6521</points>
<connection>
<GID>1504</GID>
<name>IN_3</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>302,6519,302.5,6519</points>
<connection>
<GID>1513</GID>
<name>IN_0</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>852</ID>
<shape>
<vsegment>
<ID>13</ID>
<points>234,6582.5,234,6586</points>
<connection>
<GID>1437</GID>
<name>IN_0</name></connection>
<connection>
<GID>1436</GID>
<name>SEL_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,6517,303.5,6520</points>
<intersection>6517 2</intersection>
<intersection>6520 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,6520,306,6520</points>
<connection>
<GID>1504</GID>
<name>IN_2</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,6517,303.5,6517</points>
<connection>
<GID>1514</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,6514.5,304,6519</points>
<intersection>6514.5 2</intersection>
<intersection>6519 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,6519,306,6519</points>
<connection>
<GID>1504</GID>
<name>IN_1</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,6514.5,304,6514.5</points>
<connection>
<GID>1515</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>854</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,6582.5,235,6588</points>
<connection>
<GID>1436</GID>
<name>SEL_1</name></connection>
<intersection>6588 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>234,6588,235,6588</points>
<connection>
<GID>1438</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>1244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,6512,304.5,6518</points>
<intersection>6512 2</intersection>
<intersection>6518 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,6518,306,6518</points>
<connection>
<GID>1504</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,6512,304.5,6512</points>
<connection>
<GID>1516</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>855</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,6582.5,236,6590</points>
<connection>
<GID>1436</GID>
<name>SEL_0</name></connection>
<intersection>6590 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,6590,236,6590</points>
<connection>
<GID>1439</GID>
<name>IN_0</name></connection>
<intersection>236 0</intersection></hsegment></shape></wire>
<wire>
<ID>1245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,6521.5,341.5,6521.5</points>
<connection>
<GID>1517</GID>
<name>OUT</name></connection>
<connection>
<GID>1518</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>856</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231,6570,231,6573.5</points>
<intersection>6570 2</intersection>
<intersection>6573.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>231,6573.5,232,6573.5</points>
<connection>
<GID>1436</GID>
<name>IN_0</name></connection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,6570,231,6570</points>
<connection>
<GID>1335</GID>
<name>IN_0</name></connection>
<intersection>231 0</intersection></hsegment></shape></wire>
<wire>
<ID>1246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338.5,6527,338.5,6531.5</points>
<connection>
<GID>1517</GID>
<name>SEL_1</name></connection>
<intersection>6531.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>337.5,6531.5,338.5,6531.5</points>
<connection>
<GID>1519</GID>
<name>IN_0</name></connection>
<intersection>338.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>857</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,6572,230.5,6574.5</points>
<intersection>6572 3</intersection>
<intersection>6574.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230.5,6574.5,232,6574.5</points>
<connection>
<GID>1436</GID>
<name>IN_1</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228,6572,230.5,6572</points>
<connection>
<GID>1336</GID>
<name>IN_0</name></connection>
<intersection>230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,6527,339.5,6533.5</points>
<connection>
<GID>1517</GID>
<name>SEL_0</name></connection>
<intersection>6533.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>338.5,6533.5,339.5,6533.5</points>
<connection>
<GID>1520</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>858</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,6574,230,6575.5</points>
<intersection>6574 2</intersection>
<intersection>6575.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,6575.5,232,6575.5</points>
<connection>
<GID>1436</GID>
<name>IN_2</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,6574,230,6574</points>
<connection>
<GID>1337</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>1248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,6527,337.5,6529.5</points>
<connection>
<GID>1517</GID>
<name>SEL_2</name></connection>
<intersection>6529.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336,6529.5,337.5,6529.5</points>
<connection>
<GID>1521</GID>
<name>IN_0</name></connection>
<intersection>337.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>859</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228,6576,230,6576</points>
<connection>
<GID>1338</GID>
<name>IN_0</name></connection>
<intersection>230 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>230,6576,230,6576.5</points>
<intersection>6576 1</intersection>
<intersection>6576.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>230,6576.5,232,6576.5</points>
<connection>
<GID>1436</GID>
<name>IN_3</name></connection>
<intersection>230 3</intersection></hsegment></shape></wire>
<wire>
<ID>1249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>335,6525,335.5,6525</points>
<connection>
<GID>1517</GID>
<name>IN_7</name></connection>
<intersection>335 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>335,6525,335,6527</points>
<intersection>6525 1</intersection>
<intersection>6527 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>332.5,6527,335,6527</points>
<connection>
<GID>1473</GID>
<name>IN_0</name></connection>
<intersection>335 3</intersection></hsegment></shape></wire>
<wire>
<ID>860</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231,6580.5,231,6584</points>
<intersection>6580.5 1</intersection>
<intersection>6584 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>231,6580.5,232,6580.5</points>
<connection>
<GID>1436</GID>
<name>IN_7</name></connection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,6584,231,6584</points>
<connection>
<GID>1342</GID>
<name>IN_0</name></connection>
<intersection>231 0</intersection></hsegment></shape></wire>
<wire>
<ID>1250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>331.5,6524,335.5,6524</points>
<connection>
<GID>1517</GID>
<name>IN_6</name></connection>
<intersection>331.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>331.5,6524,331.5,6525</points>
<connection>
<GID>1472</GID>
<name>IN_0</name></connection>
<intersection>6524 1</intersection></vsegment></shape></wire>
<wire>
<ID>861</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,6579.5,230.5,6582</points>
<intersection>6579.5 1</intersection>
<intersection>6582 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230.5,6579.5,232,6579.5</points>
<connection>
<GID>1436</GID>
<name>IN_6</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228,6582,230.5,6582</points>
<connection>
<GID>1341</GID>
<name>IN_0</name></connection>
<intersection>230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329.5,6523,335.5,6523</points>
<connection>
<GID>1523</GID>
<name>IN_0</name></connection>
<connection>
<GID>1517</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>862</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,6578.5,230,6580</points>
<intersection>6578.5 2</intersection>
<intersection>6580 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228,6580,230,6580</points>
<connection>
<GID>1340</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230,6578.5,232,6578.5</points>
<connection>
<GID>1436</GID>
<name>IN_5</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>1252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,6521,330,6521.5</points>
<intersection>6521 8</intersection>
<intersection>6521.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>330,6521.5,335.5,6521.5</points>
<intersection>330 0</intersection>
<intersection>335.5 9</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>330,6521,330.5,6521</points>
<connection>
<GID>1522</GID>
<name>IN_0</name></connection>
<intersection>330 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>335.5,6521.5,335.5,6522</points>
<connection>
<GID>1517</GID>
<name>IN_4</name></connection>
<intersection>6521.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>863</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228,6578,230,6578</points>
<connection>
<GID>1339</GID>
<name>IN_0</name></connection>
<intersection>230 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>230,6577.5,230,6578</points>
<intersection>6577.5 4</intersection>
<intersection>6578 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>230,6577.5,232,6577.5</points>
<connection>
<GID>1436</GID>
<name>IN_4</name></connection>
<intersection>230 3</intersection></hsegment></shape></wire>
<wire>
<ID>1253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,6519,332,6521</points>
<intersection>6519 2</intersection>
<intersection>6521 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332,6521,335.5,6521</points>
<connection>
<GID>1517</GID>
<name>IN_3</name></connection>
<intersection>332 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>331.5,6519,332,6519</points>
<connection>
<GID>1474</GID>
<name>IN_0</name></connection>
<intersection>332 0</intersection></hsegment></shape></wire>
<wire>
<ID>864</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>238,6577,239.5,6577</points>
<connection>
<GID>1436</GID>
<name>OUT</name></connection>
<connection>
<GID>1343</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,6517,333,6520</points>
<intersection>6517 2</intersection>
<intersection>6520 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,6520,335.5,6520</points>
<connection>
<GID>1517</GID>
<name>IN_2</name></connection>
<intersection>333 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330,6517,333,6517</points>
<connection>
<GID>1475</GID>
<name>IN_0</name></connection>
<intersection>333 0</intersection></hsegment></shape></wire>
<wire>
<ID>865</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>264.5,6582.5,264.5,6586</points>
<connection>
<GID>1345</GID>
<name>IN_0</name></connection>
<connection>
<GID>1344</GID>
<name>SEL_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,6514.5,333.5,6519</points>
<intersection>6514.5 2</intersection>
<intersection>6519 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333.5,6519,335.5,6519</points>
<connection>
<GID>1517</GID>
<name>IN_1</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>331,6514.5,333.5,6514.5</points>
<connection>
<GID>1476</GID>
<name>IN_0</name></connection>
<intersection>333.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>866</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,6582.5,265.5,6588</points>
<connection>
<GID>1344</GID>
<name>SEL_1</name></connection>
<intersection>6588 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>264.5,6588,265.5,6588</points>
<connection>
<GID>1346</GID>
<name>IN_0</name></connection>
<intersection>265.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,6512,334,6518</points>
<intersection>6512 2</intersection>
<intersection>6518 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334,6518,335.5,6518</points>
<connection>
<GID>1517</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330.5,6512,334,6512</points>
<connection>
<GID>1477</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>867</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,6582.5,266.5,6590</points>
<connection>
<GID>1344</GID>
<name>SEL_0</name></connection>
<intersection>6590 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,6590,266.5,6590</points>
<connection>
<GID>1347</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,6493.5,312,6493.5</points>
<connection>
<GID>1484</GID>
<name>OUT</name></connection>
<connection>
<GID>1485</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>868</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,6570,261.5,6573.5</points>
<intersection>6570 2</intersection>
<intersection>6573.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,6573.5,262.5,6573.5</points>
<connection>
<GID>1344</GID>
<name>IN_0</name></connection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>258.5,6570,261.5,6570</points>
<connection>
<GID>1348</GID>
<name>IN_0</name></connection>
<intersection>261.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,6499,309,6503.5</points>
<connection>
<GID>1484</GID>
<name>SEL_1</name></connection>
<intersection>6503.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>308,6503.5,309,6503.5</points>
<connection>
<GID>1486</GID>
<name>IN_0</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>869</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,6572,261,6574.5</points>
<intersection>6572 3</intersection>
<intersection>6574.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,6574.5,262.5,6574.5</points>
<connection>
<GID>1344</GID>
<name>IN_1</name></connection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258.5,6572,261,6572</points>
<connection>
<GID>1349</GID>
<name>IN_0</name></connection>
<intersection>261 0</intersection></hsegment></shape></wire>
<wire>
<ID>1259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,6499,310,6505.5</points>
<connection>
<GID>1484</GID>
<name>SEL_0</name></connection>
<intersection>6505.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,6505.5,310,6505.5</points>
<connection>
<GID>1487</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>870</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,6574,260.5,6575.5</points>
<intersection>6574 2</intersection>
<intersection>6575.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,6575.5,262.5,6575.5</points>
<connection>
<GID>1344</GID>
<name>IN_2</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>258.5,6574,260.5,6574</points>
<connection>
<GID>1350</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,6499,308,6501.5</points>
<connection>
<GID>1484</GID>
<name>SEL_2</name></connection>
<intersection>6501.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>306.5,6501.5,308,6501.5</points>
<connection>
<GID>1488</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>871</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258.5,6576,260.5,6576</points>
<connection>
<GID>1351</GID>
<name>IN_0</name></connection>
<intersection>260.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>260.5,6576,260.5,6576.5</points>
<intersection>6576 1</intersection>
<intersection>6576.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260.5,6576.5,262.5,6576.5</points>
<connection>
<GID>1344</GID>
<name>IN_3</name></connection>
<intersection>260.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305.5,6497,306,6497</points>
<connection>
<GID>1484</GID>
<name>IN_7</name></connection>
<intersection>305.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>305.5,6497,305.5,6499</points>
<intersection>6497 1</intersection>
<intersection>6499 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>303,6499,305.5,6499</points>
<connection>
<GID>1492</GID>
<name>IN_0</name></connection>
<intersection>305.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>872</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,6580.5,261.5,6584</points>
<intersection>6580.5 1</intersection>
<intersection>6584 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,6580.5,262.5,6580.5</points>
<connection>
<GID>1344</GID>
<name>IN_7</name></connection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>258.5,6584,261.5,6584</points>
<connection>
<GID>1355</GID>
<name>IN_0</name></connection>
<intersection>261.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>302,6496,306,6496</points>
<connection>
<GID>1484</GID>
<name>IN_6</name></connection>
<intersection>302 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>302,6496,302,6497</points>
<connection>
<GID>1491</GID>
<name>IN_0</name></connection>
<intersection>6496 1</intersection></vsegment></shape></wire>
<wire>
<ID>873</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,6579.5,261,6582</points>
<intersection>6579.5 1</intersection>
<intersection>6582 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,6579.5,262.5,6579.5</points>
<connection>
<GID>1344</GID>
<name>IN_6</name></connection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258.5,6582,261,6582</points>
<connection>
<GID>1354</GID>
<name>IN_0</name></connection>
<intersection>261 0</intersection></hsegment></shape></wire>
<wire>
<ID>1263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>300,6495,306,6495</points>
<connection>
<GID>1490</GID>
<name>IN_0</name></connection>
<connection>
<GID>1484</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>874</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,6578.5,260.5,6580</points>
<intersection>6578.5 2</intersection>
<intersection>6580 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258.5,6580,260.5,6580</points>
<connection>
<GID>1353</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>260.5,6578.5,262.5,6578.5</points>
<connection>
<GID>1344</GID>
<name>IN_5</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>300.5,6493,300.5,6493.5</points>
<intersection>6493 8</intersection>
<intersection>6493.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>300.5,6493.5,306,6493.5</points>
<intersection>300.5 0</intersection>
<intersection>306 9</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>300.5,6493,301,6493</points>
<connection>
<GID>1489</GID>
<name>IN_0</name></connection>
<intersection>300.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>306,6493.5,306,6494</points>
<connection>
<GID>1484</GID>
<name>IN_4</name></connection>
<intersection>6493.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>875</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258.5,6578,260.5,6578</points>
<connection>
<GID>1352</GID>
<name>IN_0</name></connection>
<intersection>260.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>260.5,6577.5,260.5,6578</points>
<intersection>6577.5 4</intersection>
<intersection>6578 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260.5,6577.5,262.5,6577.5</points>
<connection>
<GID>1344</GID>
<name>IN_4</name></connection>
<intersection>260.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,6491,302.5,6493</points>
<intersection>6491 4</intersection>
<intersection>6493 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,6493,306,6493</points>
<connection>
<GID>1484</GID>
<name>IN_3</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>302,6491,302.5,6491</points>
<connection>
<GID>1493</GID>
<name>IN_0</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>876</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>268.5,6577,270.5,6577</points>
<connection>
<GID>1344</GID>
<name>OUT</name></connection>
<connection>
<GID>1356</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,6489,303.5,6492</points>
<intersection>6489 2</intersection>
<intersection>6492 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,6492,306,6492</points>
<connection>
<GID>1484</GID>
<name>IN_2</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,6489,303.5,6489</points>
<connection>
<GID>1494</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>877</ID>
<shape>
<vsegment>
<ID>8</ID>
<points>233,6558.5,233,6562</points>
<connection>
<GID>1371</GID>
<name>IN_0</name></connection>
<connection>
<GID>1370</GID>
<name>SEL_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,6486.5,304,6491</points>
<intersection>6486.5 2</intersection>
<intersection>6491 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,6491,306,6491</points>
<connection>
<GID>1484</GID>
<name>IN_1</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,6486.5,304,6486.5</points>
<connection>
<GID>1495</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>1268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,6484,304.5,6490</points>
<intersection>6484 2</intersection>
<intersection>6490 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,6490,306,6490</points>
<connection>
<GID>1484</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,6484,304.5,6484</points>
<connection>
<GID>1496</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,6493.5,341.5,6493.5</points>
<connection>
<GID>1497</GID>
<name>OUT</name></connection>
<connection>
<GID>1498</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338.5,6499,338.5,6503.5</points>
<connection>
<GID>1497</GID>
<name>SEL_1</name></connection>
<intersection>6503.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>337.5,6503.5,338.5,6503.5</points>
<connection>
<GID>1499</GID>
<name>IN_0</name></connection>
<intersection>338.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,6499,339.5,6505.5</points>
<connection>
<GID>1497</GID>
<name>SEL_0</name></connection>
<intersection>6505.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>338.5,6505.5,339.5,6505.5</points>
<connection>
<GID>1500</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,6499,337.5,6501.5</points>
<connection>
<GID>1497</GID>
<name>SEL_2</name></connection>
<intersection>6501.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336,6501.5,337.5,6501.5</points>
<connection>
<GID>1501</GID>
<name>IN_0</name></connection>
<intersection>337.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>335,6497,335.5,6497</points>
<connection>
<GID>1497</GID>
<name>IN_7</name></connection>
<intersection>335 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>335,6497,335,6499</points>
<intersection>6497 1</intersection>
<intersection>6499 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>332.5,6499,335,6499</points>
<connection>
<GID>1479</GID>
<name>IN_0</name></connection>
<intersection>335 3</intersection></hsegment></shape></wire>
<wire>
<ID>1274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>331.5,6496,335.5,6496</points>
<connection>
<GID>1497</GID>
<name>IN_6</name></connection>
<intersection>331.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>331.5,6496,331.5,6497</points>
<connection>
<GID>1478</GID>
<name>IN_0</name></connection>
<intersection>6496 1</intersection></vsegment></shape></wire>
<wire>
<ID>1275</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329.5,6495,335.5,6495</points>
<connection>
<GID>1503</GID>
<name>IN_0</name></connection>
<connection>
<GID>1497</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,6493,330,6493.5</points>
<intersection>6493 8</intersection>
<intersection>6493.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>330,6493.5,335.5,6493.5</points>
<intersection>330 0</intersection>
<intersection>335.5 9</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>330,6493,330.5,6493</points>
<connection>
<GID>1502</GID>
<name>IN_0</name></connection>
<intersection>330 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>335.5,6493.5,335.5,6494</points>
<connection>
<GID>1497</GID>
<name>IN_4</name></connection>
<intersection>6493.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,6491,332,6493</points>
<intersection>6491 2</intersection>
<intersection>6493 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332,6493,335.5,6493</points>
<connection>
<GID>1497</GID>
<name>IN_3</name></connection>
<intersection>332 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>331.5,6491,332,6491</points>
<connection>
<GID>1480</GID>
<name>IN_0</name></connection>
<intersection>332 0</intersection></hsegment></shape></wire>
<wire>
<ID>1278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,6489,333,6492</points>
<intersection>6489 2</intersection>
<intersection>6492 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,6492,335.5,6492</points>
<connection>
<GID>1497</GID>
<name>IN_2</name></connection>
<intersection>333 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330,6489,333,6489</points>
<connection>
<GID>1481</GID>
<name>IN_0</name></connection>
<intersection>333 0</intersection></hsegment></shape></wire>
<wire>
<ID>1279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,6486.5,333.5,6491</points>
<intersection>6486.5 2</intersection>
<intersection>6491 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333.5,6491,335.5,6491</points>
<connection>
<GID>1497</GID>
<name>IN_1</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>331,6486.5,333.5,6486.5</points>
<connection>
<GID>1482</GID>
<name>IN_0</name></connection>
<intersection>333.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,6484,334,6490</points>
<intersection>6484 2</intersection>
<intersection>6490 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334,6490,335.5,6490</points>
<connection>
<GID>1497</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330.5,6484,334,6484</points>
<connection>
<GID>1483</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>1281</ID>
<shape>
<hsegment>
<ID>25</ID>
<points>391,6578.5,391.5,6578.5</points>
<connection>
<GID>1555</GID>
<name>IN_0</name></connection>
<connection>
<GID>1568</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1282</ID>
<shape>
<hsegment>
<ID>13</ID>
<points>391,6543.5,391.5,6543.5</points>
<connection>
<GID>1561</GID>
<name>IN_0</name></connection>
<connection>
<GID>1567</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1283</ID>
<shape>
<hsegment>
<ID>12</ID>
<points>391,6548.5,391.5,6548.5</points>
<connection>
<GID>1560</GID>
<name>IN_0</name></connection>
<connection>
<GID>1566</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1284</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>391,6553.5,391.5,6553.5</points>
<connection>
<GID>1559</GID>
<name>IN_0</name></connection>
<connection>
<GID>1565</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1285</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>391,6558.5,391.5,6558.5</points>
<connection>
<GID>1562</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1286</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>391,6563.5,391.5,6563.5</points>
<connection>
<GID>1558</GID>
<name>IN_0</name></connection>
<connection>
<GID>1563</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1287</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>391,6568.5,391.5,6568.5</points>
<connection>
<GID>1557</GID>
<name>IN_0</name></connection>
<connection>
<GID>1570</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1288</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>391,6573.5,391.5,6573.5</points>
<connection>
<GID>1556</GID>
<name>IN_0</name></connection>
<connection>
<GID>1569</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1289</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>398.5,6547,398.5,6584.5</points>
<intersection>6547 36</intersection>
<intersection>6552 44</intersection>
<intersection>6557 43</intersection>
<intersection>6562 42</intersection>
<intersection>6567 41</intersection>
<intersection>6572 40</intersection>
<intersection>6577 39</intersection>
<intersection>6582 38</intersection>
<intersection>6584.5 37</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>393.5,6547,398.5,6547</points>
<connection>
<GID>1561</GID>
<name>SEL_0</name></connection>
<intersection>398.5 3</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>393.5,6584.5,398.5,6584.5</points>
<connection>
<GID>1571</GID>
<name>IN_0</name></connection>
<intersection>398.5 3</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>393.5,6582,398.5,6582</points>
<connection>
<GID>1555</GID>
<name>SEL_0</name></connection>
<intersection>398.5 3</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>393.5,6577,398.5,6577</points>
<connection>
<GID>1556</GID>
<name>SEL_0</name></connection>
<intersection>398.5 3</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>393.5,6572,398.5,6572</points>
<connection>
<GID>1557</GID>
<name>SEL_0</name></connection>
<intersection>398.5 3</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>393.5,6567,398.5,6567</points>
<connection>
<GID>1558</GID>
<name>SEL_0</name></connection>
<intersection>398.5 3</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>393.5,6562,398.5,6562</points>
<connection>
<GID>1562</GID>
<name>SEL_0</name></connection>
<intersection>398.5 3</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>393.5,6557,398.5,6557</points>
<connection>
<GID>1559</GID>
<name>SEL_0</name></connection>
<intersection>398.5 3</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>393.5,6552,398.5,6552</points>
<connection>
<GID>1560</GID>
<name>SEL_0</name></connection>
<intersection>398.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1290</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>391,6545.5,391.5,6545.5</points>
<connection>
<GID>1561</GID>
<name>IN_1</name></connection>
<connection>
<GID>1573</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1291</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>391,6550.5,391.5,6550.5</points>
<connection>
<GID>1560</GID>
<name>IN_1</name></connection>
<connection>
<GID>1574</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1292</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>391,6555.5,391.5,6555.5</points>
<connection>
<GID>1559</GID>
<name>IN_1</name></connection>
<connection>
<GID>1575</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1293</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>391,6560.5,391.5,6560.5</points>
<connection>
<GID>1562</GID>
<name>IN_1</name></connection>
<connection>
<GID>1576</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1294</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>391,6565.5,391.5,6565.5</points>
<connection>
<GID>1558</GID>
<name>IN_1</name></connection>
<connection>
<GID>1577</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1295</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>391,6570.5,391.5,6570.5</points>
<connection>
<GID>1557</GID>
<name>IN_1</name></connection>
<connection>
<GID>1578</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1296</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>391,6575.5,391.5,6575.5</points>
<connection>
<GID>1556</GID>
<name>IN_1</name></connection>
<connection>
<GID>1579</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1297</ID>
<shape>
<hsegment>
<ID>17</ID>
<points>391,6580.5,391.5,6580.5</points>
<connection>
<GID>1555</GID>
<name>IN_1</name></connection>
<connection>
<GID>1580</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1298</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>395.5,6579.5,401.5,6579.5</points>
<connection>
<GID>1547</GID>
<name>IN_0</name></connection>
<connection>
<GID>1555</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>395.5,6574.5,401.5,6574.5</points>
<connection>
<GID>1556</GID>
<name>OUT</name></connection>
<connection>
<GID>1548</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>395.5,6569.5,401.5,6569.5</points>
<connection>
<GID>1557</GID>
<name>OUT</name></connection>
<connection>
<GID>1549</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>395.5,6564.5,401.5,6564.5</points>
<connection>
<GID>1558</GID>
<name>OUT</name></connection>
<connection>
<GID>1550</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>395.5,6559.5,401.5,6559.5</points>
<connection>
<GID>1562</GID>
<name>OUT</name></connection>
<connection>
<GID>1551</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1303</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>395.5,6554.5,401,6554.5</points>
<connection>
<GID>1559</GID>
<name>OUT</name></connection>
<connection>
<GID>1552</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1304</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>395.5,6549.5,401,6549.5</points>
<connection>
<GID>1553</GID>
<name>IN_0</name></connection>
<connection>
<GID>1560</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1305</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>395.5,6544.5,401,6544.5</points>
<connection>
<GID>1554</GID>
<name>IN_0</name></connection>
<connection>
<GID>1561</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>931</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,6558.5,234,6564</points>
<connection>
<GID>1370</GID>
<name>SEL_1</name></connection>
<intersection>6564 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>233,6564,234,6564</points>
<connection>
<GID>1372</GID>
<name>IN_0</name></connection>
<intersection>234 0</intersection></hsegment></shape></wire>
<wire>
<ID>936</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,6558.5,235,6566</points>
<connection>
<GID>1370</GID>
<name>SEL_0</name></connection>
<intersection>6566 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233,6566,235,6566</points>
<connection>
<GID>1373</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>1038</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,6546,230,6549.5</points>
<intersection>6546 2</intersection>
<intersection>6549.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,6549.5,231,6549.5</points>
<connection>
<GID>1370</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,6546,230,6546</points>
<connection>
<GID>1374</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>1039</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,6548,229.5,6550.5</points>
<intersection>6548 3</intersection>
<intersection>6550.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,6550.5,231,6550.5</points>
<connection>
<GID>1370</GID>
<name>IN_1</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>227,6548,229.5,6548</points>
<connection>
<GID>1375</GID>
<name>IN_0</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1040</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,6550,229,6551.5</points>
<intersection>6550 2</intersection>
<intersection>6551.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,6551.5,231,6551.5</points>
<connection>
<GID>1370</GID>
<name>IN_2</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,6550,229,6550</points>
<connection>
<GID>1376</GID>
<name>IN_0</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>1041</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,6552,229,6552</points>
<connection>
<GID>1377</GID>
<name>IN_0</name></connection>
<intersection>229 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229,6552,229,6552.5</points>
<intersection>6552 1</intersection>
<intersection>6552.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229,6552.5,231,6552.5</points>
<connection>
<GID>1370</GID>
<name>IN_3</name></connection>
<intersection>229 3</intersection></hsegment></shape></wire>
<wire>
<ID>1042</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,6556.5,230,6560</points>
<intersection>6556.5 1</intersection>
<intersection>6560 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,6556.5,231,6556.5</points>
<connection>
<GID>1370</GID>
<name>IN_7</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,6560,230,6560</points>
<connection>
<GID>1381</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>1043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,6555.5,229.5,6558</points>
<intersection>6555.5 1</intersection>
<intersection>6558 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,6555.5,231,6555.5</points>
<connection>
<GID>1370</GID>
<name>IN_6</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>227,6558,229.5,6558</points>
<connection>
<GID>1380</GID>
<name>IN_0</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1044</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,6554.5,229,6556</points>
<intersection>6554.5 2</intersection>
<intersection>6556 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,6556,229,6556</points>
<connection>
<GID>1379</GID>
<name>IN_0</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229,6554.5,231,6554.5</points>
<connection>
<GID>1370</GID>
<name>IN_5</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>1045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,6554,229,6554</points>
<connection>
<GID>1378</GID>
<name>IN_0</name></connection>
<intersection>229 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229,6553.5,229,6554</points>
<intersection>6553.5 4</intersection>
<intersection>6554 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229,6553.5,231,6553.5</points>
<connection>
<GID>1370</GID>
<name>IN_4</name></connection>
<intersection>229 3</intersection></hsegment></shape></wire>
<wire>
<ID>1046</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>237,6553,238.5,6553</points>
<connection>
<GID>1370</GID>
<name>OUT</name></connection>
<connection>
<GID>1382</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1047</ID>
<shape>
<vsegment>
<ID>8</ID>
<points>263.5,6558.5,263.5,6562</points>
<connection>
<GID>1358</GID>
<name>IN_0</name></connection>
<connection>
<GID>1357</GID>
<name>SEL_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1048</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,6558.5,264.5,6564</points>
<connection>
<GID>1357</GID>
<name>SEL_1</name></connection>
<intersection>6564 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>263.5,6564,264.5,6564</points>
<connection>
<GID>1359</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1049</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,6558.5,265.5,6566</points>
<connection>
<GID>1357</GID>
<name>SEL_0</name></connection>
<intersection>6566 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263.5,6566,265.5,6566</points>
<connection>
<GID>1360</GID>
<name>IN_0</name></connection>
<intersection>265.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1050</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,6546,260.5,6549.5</points>
<intersection>6546 2</intersection>
<intersection>6549.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,6549.5,261.5,6549.5</points>
<connection>
<GID>1357</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,6546,260.5,6546</points>
<connection>
<GID>1361</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1051</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,6548,260,6550.5</points>
<intersection>6548 3</intersection>
<intersection>6550.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,6550.5,261.5,6550.5</points>
<connection>
<GID>1357</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>257.5,6548,260,6548</points>
<connection>
<GID>1362</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>1052</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,6550,259.5,6551.5</points>
<intersection>6550 2</intersection>
<intersection>6551.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,6551.5,261.5,6551.5</points>
<connection>
<GID>1357</GID>
<name>IN_2</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,6550,259.5,6550</points>
<connection>
<GID>1363</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>257.5,6552,259.5,6552</points>
<connection>
<GID>1364</GID>
<name>IN_0</name></connection>
<intersection>259.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>259.5,6552,259.5,6552.5</points>
<intersection>6552 1</intersection>
<intersection>6552.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,6552.5,261.5,6552.5</points>
<connection>
<GID>1357</GID>
<name>IN_3</name></connection>
<intersection>259.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1054</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,6556.5,260.5,6560</points>
<intersection>6556.5 1</intersection>
<intersection>6560 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,6556.5,261.5,6556.5</points>
<connection>
<GID>1357</GID>
<name>IN_7</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,6560,260.5,6560</points>
<connection>
<GID>1368</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1055</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,6555.5,260,6558</points>
<intersection>6555.5 1</intersection>
<intersection>6558 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,6555.5,261.5,6555.5</points>
<connection>
<GID>1357</GID>
<name>IN_6</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>257.5,6558,260,6558</points>
<connection>
<GID>1367</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>1056</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,6554.5,259.5,6556</points>
<intersection>6554.5 2</intersection>
<intersection>6556 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,6556,259.5,6556</points>
<connection>
<GID>1366</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,6554.5,261.5,6554.5</points>
<connection>
<GID>1357</GID>
<name>IN_5</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>257.5,6554,259.5,6554</points>
<connection>
<GID>1365</GID>
<name>IN_0</name></connection>
<intersection>259.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>259.5,6553.5,259.5,6554</points>
<intersection>6553.5 4</intersection>
<intersection>6554 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,6553.5,261.5,6553.5</points>
<connection>
<GID>1357</GID>
<name>IN_4</name></connection>
<intersection>259.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1058</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>267.5,6553,269.5,6553</points>
<connection>
<GID>1357</GID>
<name>OUT</name></connection>
<connection>
<GID>1369</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1059</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>233,6534,233,6537.5</points>
<connection>
<GID>1397</GID>
<name>IN_0</name></connection>
<connection>
<GID>1396</GID>
<name>SEL_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1060</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,6534,234,6539.5</points>
<connection>
<GID>1396</GID>
<name>SEL_1</name></connection>
<intersection>6539.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>233,6539.5,234,6539.5</points>
<connection>
<GID>1398</GID>
<name>IN_0</name></connection>
<intersection>234 0</intersection></hsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,6534,235,6541.5</points>
<connection>
<GID>1396</GID>
<name>SEL_0</name></connection>
<intersection>6541.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233,6541.5,235,6541.5</points>
<connection>
<GID>1399</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,6521.5,230,6525</points>
<intersection>6521.5 2</intersection>
<intersection>6525 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,6525,231,6525</points>
<connection>
<GID>1396</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,6521.5,230,6521.5</points>
<connection>
<GID>1400</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,6523.5,229.5,6526</points>
<intersection>6523.5 3</intersection>
<intersection>6526 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,6526,231,6526</points>
<connection>
<GID>1396</GID>
<name>IN_1</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>227,6523.5,229.5,6523.5</points>
<connection>
<GID>1401</GID>
<name>IN_0</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,6525.5,229,6527</points>
<intersection>6525.5 2</intersection>
<intersection>6527 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,6527,231,6527</points>
<connection>
<GID>1396</GID>
<name>IN_2</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,6525.5,229,6525.5</points>
<connection>
<GID>1402</GID>
<name>IN_0</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,6527.5,229,6527.5</points>
<connection>
<GID>1403</GID>
<name>IN_0</name></connection>
<intersection>229 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229,6527.5,229,6528</points>
<intersection>6527.5 1</intersection>
<intersection>6528 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229,6528,231,6528</points>
<connection>
<GID>1396</GID>
<name>IN_3</name></connection>
<intersection>229 3</intersection></hsegment></shape></wire>
<wire>
<ID>1066</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,6532,230,6535.5</points>
<intersection>6532 1</intersection>
<intersection>6535.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,6532,231,6532</points>
<connection>
<GID>1396</GID>
<name>IN_7</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,6535.5,230,6535.5</points>
<connection>
<GID>1407</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>1067</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,6531,229.5,6533.5</points>
<intersection>6531 1</intersection>
<intersection>6533.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,6531,231,6531</points>
<connection>
<GID>1396</GID>
<name>IN_6</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>227,6533.5,229.5,6533.5</points>
<connection>
<GID>1406</GID>
<name>IN_0</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1068</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,6530,229,6531.5</points>
<intersection>6530 2</intersection>
<intersection>6531.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,6531.5,229,6531.5</points>
<connection>
<GID>1405</GID>
<name>IN_0</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229,6530,231,6530</points>
<connection>
<GID>1396</GID>
<name>IN_5</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>1069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,6529.5,229,6529.5</points>
<connection>
<GID>1404</GID>
<name>IN_0</name></connection>
<intersection>229 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229,6529,229,6529.5</points>
<intersection>6529 4</intersection>
<intersection>6529.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229,6529,231,6529</points>
<connection>
<GID>1396</GID>
<name>IN_4</name></connection>
<intersection>229 3</intersection></hsegment></shape></wire>
<wire>
<ID>1070</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>237,6528.5,238.5,6528.5</points>
<connection>
<GID>1396</GID>
<name>OUT</name></connection>
<connection>
<GID>1408</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1071</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>263.5,6534,263.5,6537.5</points>
<connection>
<GID>1384</GID>
<name>IN_0</name></connection>
<connection>
<GID>1383</GID>
<name>SEL_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1072</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,6534,264.5,6539.5</points>
<connection>
<GID>1383</GID>
<name>SEL_1</name></connection>
<intersection>6539.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>263.5,6539.5,264.5,6539.5</points>
<connection>
<GID>1385</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1073</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,6534,265.5,6541.5</points>
<connection>
<GID>1383</GID>
<name>SEL_0</name></connection>
<intersection>6541.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263.5,6541.5,265.5,6541.5</points>
<connection>
<GID>1386</GID>
<name>IN_0</name></connection>
<intersection>265.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1074</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,6521.5,260.5,6525</points>
<intersection>6521.5 2</intersection>
<intersection>6525 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,6525,261.5,6525</points>
<connection>
<GID>1383</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,6521.5,260.5,6521.5</points>
<connection>
<GID>1387</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1075</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,6523.5,260,6526</points>
<intersection>6523.5 3</intersection>
<intersection>6526 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,6526,261.5,6526</points>
<connection>
<GID>1383</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>257.5,6523.5,260,6523.5</points>
<connection>
<GID>1388</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>1076</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,6525.5,259.5,6527</points>
<intersection>6525.5 2</intersection>
<intersection>6527 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,6527,261.5,6527</points>
<connection>
<GID>1383</GID>
<name>IN_2</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,6525.5,259.5,6525.5</points>
<connection>
<GID>1389</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1077</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>257.5,6527.5,259.5,6527.5</points>
<connection>
<GID>1390</GID>
<name>IN_0</name></connection>
<intersection>259.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>259.5,6527.5,259.5,6528</points>
<intersection>6527.5 1</intersection>
<intersection>6528 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,6528,261.5,6528</points>
<connection>
<GID>1383</GID>
<name>IN_3</name></connection>
<intersection>259.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1078</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,6532,260.5,6535.5</points>
<intersection>6532 1</intersection>
<intersection>6535.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,6532,261.5,6532</points>
<connection>
<GID>1383</GID>
<name>IN_7</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,6535.5,260.5,6535.5</points>
<connection>
<GID>1394</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1079</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,6531,260,6533.5</points>
<intersection>6531 1</intersection>
<intersection>6533.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,6531,261.5,6531</points>
<connection>
<GID>1383</GID>
<name>IN_6</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>257.5,6533.5,260,6533.5</points>
<connection>
<GID>1393</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>1080</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,6530,259.5,6531.5</points>
<intersection>6530 2</intersection>
<intersection>6531.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,6531.5,259.5,6531.5</points>
<connection>
<GID>1392</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,6530,261.5,6530</points>
<connection>
<GID>1383</GID>
<name>IN_5</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1081</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>257.5,6529.5,259.5,6529.5</points>
<connection>
<GID>1391</GID>
<name>IN_0</name></connection>
<intersection>259.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>259.5,6529,259.5,6529.5</points>
<intersection>6529 4</intersection>
<intersection>6529.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,6529,261.5,6529</points>
<connection>
<GID>1383</GID>
<name>IN_4</name></connection>
<intersection>259.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1082</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>267.5,6528.5,269.5,6528.5</points>
<connection>
<GID>1383</GID>
<name>OUT</name></connection>
<connection>
<GID>1395</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1083</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>233,6510,233,6513.5</points>
<connection>
<GID>1423</GID>
<name>IN_0</name></connection>
<connection>
<GID>1422</GID>
<name>SEL_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1084</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,6510,234,6515.5</points>
<connection>
<GID>1422</GID>
<name>SEL_1</name></connection>
<intersection>6515.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>233,6515.5,234,6515.5</points>
<connection>
<GID>1424</GID>
<name>IN_0</name></connection>
<intersection>234 0</intersection></hsegment></shape></wire>
<wire>
<ID>1085</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,6510,235,6517.5</points>
<connection>
<GID>1422</GID>
<name>SEL_0</name></connection>
<intersection>6517.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233,6517.5,235,6517.5</points>
<connection>
<GID>1425</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>1086</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,6497.5,230,6501</points>
<intersection>6497.5 2</intersection>
<intersection>6501 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,6501,231,6501</points>
<connection>
<GID>1422</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,6497.5,230,6497.5</points>
<connection>
<GID>1426</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>1087</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,6499.5,229.5,6502</points>
<intersection>6499.5 3</intersection>
<intersection>6502 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,6502,231,6502</points>
<connection>
<GID>1422</GID>
<name>IN_1</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>227,6499.5,229.5,6499.5</points>
<connection>
<GID>1427</GID>
<name>IN_0</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1088</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,6501.5,229,6503</points>
<intersection>6501.5 2</intersection>
<intersection>6503 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,6503,231,6503</points>
<connection>
<GID>1422</GID>
<name>IN_2</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,6501.5,229,6501.5</points>
<connection>
<GID>1428</GID>
<name>IN_0</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>1089</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,6503.5,229,6503.5</points>
<connection>
<GID>1429</GID>
<name>IN_0</name></connection>
<intersection>229 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229,6503.5,229,6504</points>
<intersection>6503.5 1</intersection>
<intersection>6504 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229,6504,231,6504</points>
<connection>
<GID>1422</GID>
<name>IN_3</name></connection>
<intersection>229 3</intersection></hsegment></shape></wire>
<wire>
<ID>1090</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,6508,230,6511.5</points>
<intersection>6508 1</intersection>
<intersection>6511.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,6508,231,6508</points>
<connection>
<GID>1422</GID>
<name>IN_7</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,6511.5,230,6511.5</points>
<connection>
<GID>1433</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>1091</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,6507,229.5,6509.5</points>
<intersection>6507 1</intersection>
<intersection>6509.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,6507,231,6507</points>
<connection>
<GID>1422</GID>
<name>IN_6</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>227,6509.5,229.5,6509.5</points>
<connection>
<GID>1432</GID>
<name>IN_0</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1092</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,6506,229,6507.5</points>
<intersection>6506 2</intersection>
<intersection>6507.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,6507.5,229,6507.5</points>
<connection>
<GID>1431</GID>
<name>IN_0</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229,6506,231,6506</points>
<connection>
<GID>1422</GID>
<name>IN_5</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>1093</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,6505.5,229,6505.5</points>
<connection>
<GID>1430</GID>
<name>IN_0</name></connection>
<intersection>229 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229,6505,229,6505.5</points>
<intersection>6505 4</intersection>
<intersection>6505.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229,6505,231,6505</points>
<connection>
<GID>1422</GID>
<name>IN_4</name></connection>
<intersection>229 3</intersection></hsegment></shape></wire>
<wire>
<ID>1094</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>237,6504.5,238.5,6504.5</points>
<connection>
<GID>1422</GID>
<name>OUT</name></connection>
<connection>
<GID>1434</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1095</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>263.5,6510,263.5,6513.5</points>
<connection>
<GID>1410</GID>
<name>IN_0</name></connection>
<connection>
<GID>1409</GID>
<name>SEL_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1096</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,6510,264.5,6515.5</points>
<connection>
<GID>1409</GID>
<name>SEL_1</name></connection>
<intersection>6515.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>263.5,6515.5,264.5,6515.5</points>
<connection>
<GID>1411</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1097</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>388.5,6493,392.5,6493</points>
<connection>
<GID>1240</GID>
<name>IN_0</name></connection>
<connection>
<GID>1242</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1098</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,6510,265.5,6517.5</points>
<connection>
<GID>1409</GID>
<name>SEL_0</name></connection>
<intersection>6517.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263.5,6517.5,265.5,6517.5</points>
<connection>
<GID>1412</GID>
<name>IN_0</name></connection>
<intersection>265.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1099</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>400,6509,401.5,6509</points>
<connection>
<GID>1225</GID>
<name>OUT</name></connection>
<connection>
<GID>1227</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1100</ID>
<shape>
<hsegment>
<ID>21</ID>
<points>427.5,6513.5,428.5,6513.5</points>
<connection>
<GID>1215</GID>
<name>OUT</name></connection>
<connection>
<GID>1228</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>417,6506.5,417,6510</points>
<intersection>6506.5 1</intersection>
<intersection>6510 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>413,6506.5,417,6506.5</points>
<connection>
<GID>1223</GID>
<name>IN_0</name></connection>
<intersection>417 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>417,6510,420.5,6510</points>
<connection>
<GID>1215</GID>
<name>IN_4</name></connection>
<intersection>417 0</intersection></hsegment></shape></wire>
<wire>
<ID>1102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>392,6504.5,392,6506.5</points>
<intersection>6504.5 3</intersection>
<intersection>6506.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>392,6506.5,394,6506.5</points>
<connection>
<GID>1225</GID>
<name>IN_1</name></connection>
<intersection>392 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>388.5,6504.5,392,6504.5</points>
<connection>
<GID>1230</GID>
<name>IN_0</name></connection>
<intersection>392 0</intersection></hsegment></shape></wire>
<wire>
<ID>1103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>391,6507.5,394,6507.5</points>
<connection>
<GID>1225</GID>
<name>IN_2</name></connection>
<intersection>391 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>391,6506.5,391,6507.5</points>
<intersection>6506.5 6</intersection>
<intersection>6507.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>388.5,6506.5,391,6506.5</points>
<connection>
<GID>1231</GID>
<name>IN_0</name></connection>
<intersection>391 5</intersection></hsegment></shape></wire>
<wire>
<ID>1104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>388.5,6508.5,394,6508.5</points>
<connection>
<GID>1225</GID>
<name>IN_3</name></connection>
<connection>
<GID>1229</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>388.5,6510.5,394,6510.5</points>
<connection>
<GID>1225</GID>
<name>IN_5</name></connection>
<connection>
<GID>1233</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>391,6511.5,394,6511.5</points>
<connection>
<GID>1225</GID>
<name>IN_6</name></connection>
<intersection>391 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>391,6511.5,391,6512.5</points>
<intersection>6511.5 1</intersection>
<intersection>6512.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>388.5,6512.5,391,6512.5</points>
<connection>
<GID>1232</GID>
<name>IN_0</name></connection>
<intersection>391 4</intersection></hsegment></shape></wire>
<wire>
<ID>1107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>392,6512.5,392,6514.5</points>
<intersection>6512.5 1</intersection>
<intersection>6514.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>392,6512.5,394,6512.5</points>
<connection>
<GID>1225</GID>
<name>IN_7</name></connection>
<intersection>392 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>388.5,6514.5,392,6514.5</points>
<connection>
<GID>1234</GID>
<name>IN_0</name></connection>
<intersection>392 0</intersection></hsegment></shape></wire>
<wire>
<ID>1108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>395,6517,396,6517</points>
<connection>
<GID>1236</GID>
<name>IN_0</name></connection>
<intersection>396 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>396,6514.5,396,6517</points>
<connection>
<GID>1225</GID>
<name>SEL_2</name></connection>
<intersection>6517 1</intersection></vsegment></shape></wire>
<wire>
<ID>1109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397,6514.5,397,6519</points>
<connection>
<GID>1225</GID>
<name>SEL_1</name></connection>
<intersection>6519 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>395,6519,397,6519</points>
<connection>
<GID>1237</GID>
<name>IN_0</name></connection>
<intersection>397 0</intersection></hsegment></shape></wire>
<wire>
<ID>1110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,6514.5,398,6521</points>
<connection>
<GID>1225</GID>
<name>SEL_0</name></connection>
<intersection>6521 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>395,6521,398,6521</points>
<connection>
<GID>1235</GID>
<name>IN_0</name></connection>
<intersection>398 0</intersection></hsegment></shape></wire>
<wire>
<ID>1111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>390,6503,390,6509.5</points>
<connection>
<GID>1238</GID>
<name>OUT_0</name></connection>
<intersection>6505.5 6</intersection>
<intersection>6509.5 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>390,6505.5,394,6505.5</points>
<connection>
<GID>1225</GID>
<name>IN_0</name></connection>
<intersection>390 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>390,6509.5,394,6509.5</points>
<connection>
<GID>1225</GID>
<name>IN_4</name></connection>
<intersection>390 0</intersection></hsegment></shape></wire>
<wire>
<ID>1112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>419.5,6489.5,419.5,6492</points>
<intersection>6489.5 5</intersection>
<intersection>6492 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>419.5,6492,421,6492</points>
<connection>
<GID>1239</GID>
<name>IN_1</name></connection>
<intersection>419.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>418.5,6489.5,419.5,6489.5</points>
<connection>
<GID>1241</GID>
<name>OUT</name></connection>
<intersection>419.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1113</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>410,6497.5,410,6498.5</points>
<intersection>6497.5 11</intersection>
<intersection>6498.5 12</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>410,6497.5,412.5,6497.5</points>
<connection>
<GID>1243</GID>
<name>IN_0</name></connection>
<intersection>410 10</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>408.5,6498.5,410,6498.5</points>
<connection>
<GID>1244</GID>
<name>IN_0</name></connection>
<intersection>410 10</intersection></hsegment></shape></wire>
<wire>
<ID>1114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>419.5,6494,421,6494</points>
<connection>
<GID>1239</GID>
<name>IN_0</name></connection>
<intersection>419.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>419.5,6494,419.5,6496.5</points>
<intersection>6494 1</intersection>
<intersection>6496.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>418.5,6496.5,419.5,6496.5</points>
<connection>
<GID>1243</GID>
<name>OUT</name></connection>
<intersection>419.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410,6490.5,412.5,6490.5</points>
<connection>
<GID>1241</GID>
<name>IN_0</name></connection>
<intersection>410 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>410,6490.5,410,6491</points>
<intersection>6490.5 1</intersection>
<intersection>6491 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>408.5,6491,410,6491</points>
<connection>
<GID>1245</GID>
<name>IN_0</name></connection>
<intersection>410 12</intersection></hsegment></shape></wire>
<wire>
<ID>1116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>410,6494.5,410,6495.5</points>
<intersection>6494.5 3</intersection>
<intersection>6495.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>410,6495.5,412.5,6495.5</points>
<connection>
<GID>1243</GID>
<name>IN_1</name></connection>
<intersection>410 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>408.5,6494.5,410,6494.5</points>
<connection>
<GID>1246</GID>
<name>IN_0</name></connection>
<intersection>410 0</intersection></hsegment></shape></wire>
<wire>
<ID>1117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410,6488.5,412.5,6488.5</points>
<connection>
<GID>1241</GID>
<name>IN_1</name></connection>
<intersection>410 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>410,6488,410,6488.5</points>
<intersection>6488 6</intersection>
<intersection>6488.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>408.5,6488,410,6488</points>
<connection>
<GID>1247</GID>
<name>IN_0</name></connection>
<intersection>410 4</intersection></hsegment></shape></wire>
<wire>
<ID>1118</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>427,6493,428.5,6493</points>
<connection>
<GID>1239</GID>
<name>OUT</name></connection>
<connection>
<GID>1248</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>413,6520.5,417,6520.5</points>
<connection>
<GID>1216</GID>
<name>IN_0</name></connection>
<intersection>417 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>417,6517,417,6520.5</points>
<intersection>6517 4</intersection>
<intersection>6520.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>417,6517,420.5,6517</points>
<connection>
<GID>1215</GID>
<name>IN_0</name></connection>
<intersection>417 3</intersection></hsegment></shape></wire>
<wire>
<ID>1120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>416.5,6508.5,416.5,6511</points>
<intersection>6508.5 3</intersection>
<intersection>6511 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>416.5,6511,420.5,6511</points>
<connection>
<GID>1215</GID>
<name>IN_5</name></connection>
<intersection>416.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>413,6508.5,416.5,6508.5</points>
<connection>
<GID>1222</GID>
<name>IN_0</name></connection>
<intersection>416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>416,6510.5,416,6512</points>
<intersection>6510.5 1</intersection>
<intersection>6512 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>413,6510.5,416,6510.5</points>
<connection>
<GID>1219</GID>
<name>IN_0</name></connection>
<intersection>416 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>416,6512,420.5,6512</points>
<connection>
<GID>1215</GID>
<name>IN_6</name></connection>
<intersection>416 0</intersection></hsegment></shape></wire>
<wire>
<ID>1122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>416.5,6516,416.5,6518.5</points>
<intersection>6516 2</intersection>
<intersection>6518.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>416.5,6516,420.5,6516</points>
<connection>
<GID>1215</GID>
<name>IN_1</name></connection>
<intersection>416.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>413,6518.5,416.5,6518.5</points>
<connection>
<GID>1217</GID>
<name>IN_0</name></connection>
<intersection>416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>416,6515,416,6516.5</points>
<intersection>6515 2</intersection>
<intersection>6516.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>413,6516.5,416,6516.5</points>
<connection>
<GID>1221</GID>
<name>IN_0</name></connection>
<intersection>416 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>416,6515,420.5,6515</points>
<connection>
<GID>1215</GID>
<name>IN_2</name></connection>
<intersection>416 0</intersection></hsegment></shape></wire>
<wire>
<ID>1124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415.5,6514,420.5,6514</points>
<connection>
<GID>1215</GID>
<name>IN_3</name></connection>
<intersection>415.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>415.5,6514,415.5,6514.5</points>
<intersection>6514 1</intersection>
<intersection>6514.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>413,6514.5,415.5,6514.5</points>
<connection>
<GID>1218</GID>
<name>IN_0</name></connection>
<intersection>415.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>1125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>413,6512.5,415.5,6512.5</points>
<connection>
<GID>1220</GID>
<name>IN_0</name></connection>
<intersection>415.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>415.5,6512.5,415.5,6513</points>
<intersection>6512.5 1</intersection>
<intersection>6513 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>415.5,6513,420.5,6513</points>
<connection>
<GID>1215</GID>
<name>IN_7</name></connection>
<intersection>415.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,6497.5,260.5,6501</points>
<intersection>6497.5 2</intersection>
<intersection>6501 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,6501,261.5,6501</points>
<connection>
<GID>1409</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,6497.5,260.5,6497.5</points>
<connection>
<GID>1413</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,6499.5,260,6502</points>
<intersection>6499.5 3</intersection>
<intersection>6502 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,6502,261.5,6502</points>
<connection>
<GID>1409</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>257.5,6499.5,260,6499.5</points>
<connection>
<GID>1414</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-12.9721,556.521,1765.03,-352.479</PageViewport></page 4>
<page 5>
<PageViewport>-0.25,0.275735,14.5667,-7.29926</PageViewport></page 5>
<page 6>
<PageViewport>-36.5709,10474.7,1741.43,9565.72</PageViewport></page 6>
<page 7>
<PageViewport>-36.5709,10474.7,1741.43,9565.72</PageViewport></page 7>
<page 8>
<PageViewport>-36.5709,10474.7,1741.43,9565.72</PageViewport></page 8>
<page 9>
<PageViewport>-36.5709,10474.7,1741.43,9565.72</PageViewport></page 9></circuit>